VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO D2DAdapter
  CLASS BLOCK ;
  FOREIGN D2DAdapter ;
  ORIGIN 0.000 0.000 ;
  SIZE 1314.840 BY 1325.560 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 10.640 947.540 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 10.640 1101.140 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.140 10.640 1254.740 1314.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 1309.400 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 1309.400 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 1309.400 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 1309.400 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 1309.400 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 795.930 1309.400 797.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 949.110 1309.400 950.710 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1102.290 1309.400 1103.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1255.470 1309.400 1257.070 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1314.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 1309.400 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 1309.400 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 1309.400 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 1309.400 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 1309.400 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 792.630 1309.400 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 945.810 1309.400 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1098.990 1309.400 1100.590 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1252.170 1309.400 1253.770 ;
    END
  END VPWR
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1.000 963.150 4.000 ;
    END
  END clock
  PIN io_fdi_lpClkAck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 431.840 4.000 432.440 ;
    END
  END io_fdi_lpClkAck
  PIN io_fdi_lpConfigCredit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 319.640 1313.840 320.240 ;
    END
  END io_fdi_lpConfigCredit
  PIN io_fdi_lpConfig_bits[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 278.840 1313.840 279.440 ;
    END
  END io_fdi_lpConfig_bits[0]
  PIN io_fdi_lpConfig_bits[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 788.840 4.000 789.440 ;
    END
  END io_fdi_lpConfig_bits[10]
  PIN io_fdi_lpConfig_bits[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 1321.560 734.530 1324.560 ;
    END
  END io_fdi_lpConfig_bits[11]
  PIN io_fdi_lpConfig_bits[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1.000 625.050 4.000 ;
    END
  END io_fdi_lpConfig_bits[12]
  PIN io_fdi_lpConfig_bits[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1321.560 744.190 1324.560 ;
    END
  END io_fdi_lpConfig_bits[13]
  PIN io_fdi_lpConfig_bits[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1.000 798.930 4.000 ;
    END
  END io_fdi_lpConfig_bits[14]
  PIN io_fdi_lpConfig_bits[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 387.640 4.000 388.240 ;
    END
  END io_fdi_lpConfig_bits[15]
  PIN io_fdi_lpConfig_bits[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1.000 1169.230 4.000 ;
    END
  END io_fdi_lpConfig_bits[16]
  PIN io_fdi_lpConfig_bits[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 159.840 1313.840 160.440 ;
    END
  END io_fdi_lpConfig_bits[17]
  PIN io_fdi_lpConfig_bits[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 1321.560 396.430 1324.560 ;
    END
  END io_fdi_lpConfig_bits[18]
  PIN io_fdi_lpConfig_bits[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1321.560 879.430 1324.560 ;
    END
  END io_fdi_lpConfig_bits[19]
  PIN io_fdi_lpConfig_bits[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 720.840 1313.840 721.440 ;
    END
  END io_fdi_lpConfig_bits[1]
  PIN io_fdi_lpConfig_bits[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 200.640 1313.840 201.240 ;
    END
  END io_fdi_lpConfig_bits[20]
  PIN io_fdi_lpConfig_bits[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 173.440 4.000 174.040 ;
    END
  END io_fdi_lpConfig_bits[21]
  PIN io_fdi_lpConfig_bits[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1.000 943.830 4.000 ;
    END
  END io_fdi_lpConfig_bits[22]
  PIN io_fdi_lpConfig_bits[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 812.640 4.000 813.240 ;
    END
  END io_fdi_lpConfig_bits[23]
  PIN io_fdi_lpConfig_bits[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 1.000 901.970 4.000 ;
    END
  END io_fdi_lpConfig_bits[24]
  PIN io_fdi_lpConfig_bits[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 149.640 4.000 150.240 ;
    END
  END io_fdi_lpConfig_bits[25]
  PIN io_fdi_lpConfig_bits[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1.000 367.450 4.000 ;
    END
  END io_fdi_lpConfig_bits[26]
  PIN io_fdi_lpConfig_bits[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1.000 39.010 4.000 ;
    END
  END io_fdi_lpConfig_bits[27]
  PIN io_fdi_lpConfig_bits[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1321.560 171.030 1324.560 ;
    END
  END io_fdi_lpConfig_bits[28]
  PIN io_fdi_lpConfig_bits[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1321.560 518.790 1324.560 ;
    END
  END io_fdi_lpConfig_bits[29]
  PIN io_fdi_lpConfig_bits[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1.000 1108.050 4.000 ;
    END
  END io_fdi_lpConfig_bits[2]
  PIN io_fdi_lpConfig_bits[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 268.640 4.000 269.240 ;
    END
  END io_fdi_lpConfig_bits[30]
  PIN io_fdi_lpConfig_bits[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 81.640 1313.840 82.240 ;
    END
  END io_fdi_lpConfig_bits[31]
  PIN io_fdi_lpConfig_bits[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1298.840 4.000 1299.440 ;
    END
  END io_fdi_lpConfig_bits[3]
  PIN io_fdi_lpConfig_bits[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 601.840 1313.840 602.440 ;
    END
  END io_fdi_lpConfig_bits[4]
  PIN io_fdi_lpConfig_bits[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1.000 460.830 4.000 ;
    END
  END io_fdi_lpConfig_bits[5]
  PIN io_fdi_lpConfig_bits[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1321.560 1217.530 1324.560 ;
    END
  END io_fdi_lpConfig_bits[6]
  PIN io_fdi_lpConfig_bits[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1176.440 1313.840 1177.040 ;
    END
  END io_fdi_lpConfig_bits[7]
  PIN io_fdi_lpConfig_bits[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 1321.560 1156.350 1324.560 ;
    END
  END io_fdi_lpConfig_bits[8]
  PIN io_fdi_lpConfig_bits[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1268.240 4.000 1268.840 ;
    END
  END io_fdi_lpConfig_bits[9]
  PIN io_fdi_lpConfig_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1.000 380.330 4.000 ;
    END
  END io_fdi_lpConfig_valid
  PIN io_fdi_lpCorruptCrc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 537.240 1313.840 537.840 ;
    END
  END io_fdi_lpCorruptCrc
  PIN io_fdi_lpData_bits[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1.000 1201.430 4.000 ;
    END
  END io_fdi_lpData_bits[0]
  PIN io_fdi_lpData_bits[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 452.240 1313.840 452.840 ;
    END
  END io_fdi_lpData_bits[10]
  PIN io_fdi_lpData_bits[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 1321.560 724.870 1324.560 ;
    END
  END io_fdi_lpData_bits[11]
  PIN io_fdi_lpData_bits[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1321.560 631.490 1324.560 ;
    END
  END io_fdi_lpData_bits[12]
  PIN io_fdi_lpData_bits[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 1321.560 1310.910 1324.560 ;
    END
  END io_fdi_lpData_bits[13]
  PIN io_fdi_lpData_bits[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1321.560 148.490 1324.560 ;
    END
  END io_fdi_lpData_bits[14]
  PIN io_fdi_lpData_bits[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1111.840 1313.840 1112.440 ;
    END
  END io_fdi_lpData_bits[15]
  PIN io_fdi_lpData_bits[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1321.560 35.790 1324.560 ;
    END
  END io_fdi_lpData_bits[16]
  PIN io_fdi_lpData_bits[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 615.440 1313.840 616.040 ;
    END
  END io_fdi_lpData_bits[17]
  PIN io_fdi_lpData_bits[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1.000 605.730 4.000 ;
    END
  END io_fdi_lpData_bits[18]
  PIN io_fdi_lpData_bits[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 690.240 1313.840 690.840 ;
    END
  END io_fdi_lpData_bits[19]
  PIN io_fdi_lpData_bits[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1156.040 1313.840 1156.640 ;
    END
  END io_fdi_lpData_bits[1]
  PIN io_fdi_lpData_bits[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1.000 1252.950 4.000 ;
    END
  END io_fdi_lpData_bits[20]
  PIN io_fdi_lpData_bits[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 1.000 686.230 4.000 ;
    END
  END io_fdi_lpData_bits[21]
  PIN io_fdi_lpData_bits[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 170.040 1313.840 170.640 ;
    END
  END io_fdi_lpData_bits[22]
  PIN io_fdi_lpData_bits[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 962.240 1313.840 962.840 ;
    END
  END io_fdi_lpData_bits[23]
  PIN io_fdi_lpData_bits[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1321.560 87.310 1324.560 ;
    END
  END io_fdi_lpData_bits[24]
  PIN io_fdi_lpData_bits[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 639.240 4.000 639.840 ;
    END
  END io_fdi_lpData_bits[25]
  PIN io_fdi_lpData_bits[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 584.840 4.000 585.440 ;
    END
  END io_fdi_lpData_bits[26]
  PIN io_fdi_lpData_bits[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1321.560 241.870 1324.560 ;
    END
  END io_fdi_lpData_bits[27]
  PIN io_fdi_lpData_bits[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1105.040 4.000 1105.640 ;
    END
  END io_fdi_lpData_bits[28]
  PIN io_fdi_lpData_bits[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1321.560 550.990 1324.560 ;
    END
  END io_fdi_lpData_bits[29]
  PIN io_fdi_lpData_bits[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1.000 183.910 4.000 ;
    END
  END io_fdi_lpData_bits[2]
  PIN io_fdi_lpData_bits[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 758.240 4.000 758.840 ;
    END
  END io_fdi_lpData_bits[30]
  PIN io_fdi_lpData_bits[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 1.000 1220.750 4.000 ;
    END
  END io_fdi_lpData_bits[31]
  PIN io_fdi_lpData_bits[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 1.000 995.350 4.000 ;
    END
  END io_fdi_lpData_bits[32]
  PIN io_fdi_lpData_bits[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 754.840 1313.840 755.440 ;
    END
  END io_fdi_lpData_bits[33]
  PIN io_fdi_lpData_bits[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1321.560 480.150 1324.560 ;
    END
  END io_fdi_lpData_bits[34]
  PIN io_fdi_lpData_bits[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 1.000 245.090 4.000 ;
    END
  END io_fdi_lpData_bits[35]
  PIN io_fdi_lpData_bits[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 119.040 4.000 119.640 ;
    END
  END io_fdi_lpData_bits[36]
  PIN io_fdi_lpData_bits[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 20.440 4.000 21.040 ;
    END
  END io_fdi_lpData_bits[37]
  PIN io_fdi_lpData_bits[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 204.040 4.000 204.640 ;
    END
  END io_fdi_lpData_bits[38]
  PIN io_fdi_lpData_bits[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 343.440 1313.840 344.040 ;
    END
  END io_fdi_lpData_bits[39]
  PIN io_fdi_lpData_bits[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1101.640 1313.840 1102.240 ;
    END
  END io_fdi_lpData_bits[3]
  PIN io_fdi_lpData_bits[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 1321.560 1043.650 1324.560 ;
    END
  END io_fdi_lpData_bits[40]
  PIN io_fdi_lpData_bits[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 877.240 4.000 877.840 ;
    END
  END io_fdi_lpData_bits[41]
  PIN io_fdi_lpData_bits[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1285.240 1313.840 1285.840 ;
    END
  END io_fdi_lpData_bits[42]
  PIN io_fdi_lpData_bits[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1.000 164.590 4.000 ;
    END
  END io_fdi_lpData_bits[43]
  PIN io_fdi_lpData_bits[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 693.640 4.000 694.240 ;
    END
  END io_fdi_lpData_bits[44]
  PIN io_fdi_lpData_bits[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1060.840 4.000 1061.440 ;
    END
  END io_fdi_lpData_bits[45]
  PIN io_fdi_lpData_bits[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 40.840 1313.840 41.440 ;
    END
  END io_fdi_lpData_bits[46]
  PIN io_fdi_lpData_bits[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1321.560 1001.790 1324.560 ;
    END
  END io_fdi_lpData_bits[47]
  PIN io_fdi_lpData_bits[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 1321.560 889.090 1324.560 ;
    END
  END io_fdi_lpData_bits[48]
  PIN io_fdi_lpData_bits[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 452.240 4.000 452.840 ;
    END
  END io_fdi_lpData_bits[49]
  PIN io_fdi_lpData_bits[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 442.040 1313.840 442.640 ;
    END
  END io_fdi_lpData_bits[4]
  PIN io_fdi_lpData_bits[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 1.000 132.390 4.000 ;
    END
  END io_fdi_lpData_bits[50]
  PIN io_fdi_lpData_bits[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1.000 235.430 4.000 ;
    END
  END io_fdi_lpData_bits[51]
  PIN io_fdi_lpData_bits[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 1.000 1037.210 4.000 ;
    END
  END io_fdi_lpData_bits[52]
  PIN io_fdi_lpData_bits[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 1.000 850.450 4.000 ;
    END
  END io_fdi_lpData_bits[53]
  PIN io_fdi_lpData_bits[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 496.440 4.000 497.040 ;
    END
  END io_fdi_lpData_bits[54]
  PIN io_fdi_lpData_bits[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 1.000 840.790 4.000 ;
    END
  END io_fdi_lpData_bits[55]
  PIN io_fdi_lpData_bits[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1321.560 808.590 1324.560 ;
    END
  END io_fdi_lpData_bits[56]
  PIN io_fdi_lpData_bits[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1321.560 757.070 1324.560 ;
    END
  END io_fdi_lpData_bits[57]
  PIN io_fdi_lpData_bits[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1321.560 274.070 1324.560 ;
    END
  END io_fdi_lpData_bits[58]
  PIN io_fdi_lpData_bits[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 938.440 1313.840 939.040 ;
    END
  END io_fdi_lpData_bits[59]
  PIN io_fdi_lpData_bits[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1321.560 570.310 1324.560 ;
    END
  END io_fdi_lpData_bits[5]
  PIN io_fdi_lpData_bits[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1.000 634.710 4.000 ;
    END
  END io_fdi_lpData_bits[60]
  PIN io_fdi_lpData_bits[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 1.000 1014.670 4.000 ;
    END
  END io_fdi_lpData_bits[61]
  PIN io_fdi_lpData_bits[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 180.240 1313.840 180.840 ;
    END
  END io_fdi_lpData_bits[62]
  PIN io_fdi_lpData_bits[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 105.440 1313.840 106.040 ;
    END
  END io_fdi_lpData_bits[63]
  PIN io_fdi_lpData_bits[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 1321.560 1075.850 1324.560 ;
    END
  END io_fdi_lpData_bits[6]
  PIN io_fdi_lpData_bits[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1.000 80.870 4.000 ;
    END
  END io_fdi_lpData_bits[7]
  PIN io_fdi_lpData_bits[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 418.240 1313.840 418.840 ;
    END
  END io_fdi_lpData_bits[8]
  PIN io_fdi_lpData_bits[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 928.240 1313.840 928.840 ;
    END
  END io_fdi_lpData_bits[9]
  PIN io_fdi_lpData_irdy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1200.240 1313.840 1200.840 ;
    END
  END io_fdi_lpData_irdy
  PIN io_fdi_lpData_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1149.240 4.000 1149.840 ;
    END
  END io_fdi_lpData_ready
  PIN io_fdi_lpData_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1.000 428.630 4.000 ;
    END
  END io_fdi_lpData_valid
  PIN io_fdi_lpDllpOfc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 248.240 4.000 248.840 ;
    END
  END io_fdi_lpDllpOfc
  PIN io_fdi_lpDllp_bits[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 1.000 924.510 4.000 ;
    END
  END io_fdi_lpDllp_bits[0]
  PIN io_fdi_lpDllp_bits[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 224.440 1313.840 225.040 ;
    END
  END io_fdi_lpDllp_bits[1]
  PIN io_fdi_lpDllp_bits[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1321.560 77.650 1324.560 ;
    END
  END io_fdi_lpDllp_bits[2]
  PIN io_fdi_lpDllp_bits[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1179.840 4.000 1180.440 ;
    END
  END io_fdi_lpDllp_bits[3]
  PIN io_fdi_lpDllp_bits[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 1.000 789.270 4.000 ;
    END
  END io_fdi_lpDllp_bits[4]
  PIN io_fdi_lpDllp_bits[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 309.440 1313.840 310.040 ;
    END
  END io_fdi_lpDllp_bits[5]
  PIN io_fdi_lpDllp_bits[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1321.560 860.110 1324.560 ;
    END
  END io_fdi_lpDllp_bits[6]
  PIN io_fdi_lpDllp_bits[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 258.440 4.000 259.040 ;
    END
  END io_fdi_lpDllp_bits[7]
  PIN io_fdi_lpDllp_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 442.040 4.000 442.640 ;
    END
  END io_fdi_lpDllp_valid
  PIN io_fdi_lpLinkError
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 833.040 4.000 833.640 ;
    END
  END io_fdi_lpLinkError
  PIN io_fdi_lpRetimerCrd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 115.640 1313.840 116.240 ;
    END
  END io_fdi_lpRetimerCrd
  PIN io_fdi_lpRxActiveStatus
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 1.000 1314.130 4.000 ;
    END
  END io_fdi_lpRxActiveStatus
  PIN io_fdi_lpStallAck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 646.040 1313.840 646.640 ;
    END
  END io_fdi_lpStallAck
  PIN io_fdi_lpStateReq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 680.040 1313.840 680.640 ;
    END
  END io_fdi_lpStateReq[0]
  PIN io_fdi_lpStateReq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 778.640 4.000 779.240 ;
    END
  END io_fdi_lpStateReq[1]
  PIN io_fdi_lpStateReq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1.000 113.070 4.000 ;
    END
  END io_fdi_lpStateReq[2]
  PIN io_fdi_lpStateReq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1.000 1240.070 4.000 ;
    END
  END io_fdi_lpStateReq[3]
  PIN io_fdi_lpStream_protoStack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 1.000 296.610 4.000 ;
    END
  END io_fdi_lpStream_protoStack
  PIN io_fdi_lpStream_protoType[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1321.560 786.050 1324.560 ;
    END
  END io_fdi_lpStream_protoType[0]
  PIN io_fdi_lpStream_protoType[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 561.040 1313.840 561.640 ;
    END
  END io_fdi_lpStream_protoType[1]
  PIN io_fdi_lpStream_protoType[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 1321.560 972.810 1324.560 ;
    END
  END io_fdi_lpStream_protoType[2]
  PIN io_fdi_lpWakeReq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 527.040 1313.840 527.640 ;
    END
  END io_fdi_lpWakeReq
  PIN io_fdi_plCerror
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 1.000 1281.930 4.000 ;
    END
  END io_fdi_plCerror
  PIN io_fdi_plClkReq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1321.560 222.550 1324.560 ;
    END
  END io_fdi_plClkReq
  PIN io_fdi_plConfigCredit
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1.000 225.770 4.000 ;
    END
  END io_fdi_plConfigCredit
  PIN io_fdi_plConfig_bits[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1321.560 528.450 1324.560 ;
    END
  END io_fdi_plConfig_bits[0]
  PIN io_fdi_plConfig_bits[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1.000 306.270 4.000 ;
    END
  END io_fdi_plConfig_bits[10]
  PIN io_fdi_plConfig_bits[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1094.840 4.000 1095.440 ;
    END
  END io_fdi_plConfig_bits[11]
  PIN io_fdi_plConfig_bits[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 493.040 1313.840 493.640 ;
    END
  END io_fdi_plConfig_bits[12]
  PIN io_fdi_plConfig_bits[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1321.560 654.030 1324.560 ;
    END
  END io_fdi_plConfig_bits[13]
  PIN io_fdi_plConfig_bits[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1.000 747.410 4.000 ;
    END
  END io_fdi_plConfig_bits[14]
  PIN io_fdi_plConfig_bits[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1321.560 940.610 1324.560 ;
    END
  END io_fdi_plConfig_bits[15]
  PIN io_fdi_plConfig_bits[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 734.440 1313.840 735.040 ;
    END
  END io_fdi_plConfig_bits[16]
  PIN io_fdi_plConfig_bits[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 986.040 4.000 986.640 ;
    END
  END io_fdi_plConfig_bits[17]
  PIN io_fdi_plConfig_bits[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 649.440 4.000 650.040 ;
    END
  END io_fdi_plConfig_bits[18]
  PIN io_fdi_plConfig_bits[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 129.240 4.000 129.840 ;
    END
  END io_fdi_plConfig_bits[19]
  PIN io_fdi_plConfig_bits[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1321.560 1024.330 1324.560 ;
    END
  END io_fdi_plConfig_bits[1]
  PIN io_fdi_plConfig_bits[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1.000 193.570 4.000 ;
    END
  END io_fdi_plConfig_bits[20]
  PIN io_fdi_plConfig_bits[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 1.000 1230.410 4.000 ;
    END
  END io_fdi_plConfig_bits[21]
  PIN io_fdi_plConfig_bits[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 71.440 1313.840 72.040 ;
    END
  END io_fdi_plConfig_bits[22]
  PIN io_fdi_plConfig_bits[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 64.640 4.000 65.240 ;
    END
  END io_fdi_plConfig_bits[23]
  PIN io_fdi_plConfig_bits[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 799.040 1313.840 799.640 ;
    END
  END io_fdi_plConfig_bits[24]
  PIN io_fdi_plConfig_bits[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1322.640 4.000 1323.240 ;
    END
  END io_fdi_plConfig_bits[25]
  PIN io_fdi_plConfig_bits[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1278.440 4.000 1279.040 ;
    END
  END io_fdi_plConfig_bits[26]
  PIN io_fdi_plConfig_bits[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 1321.560 1198.210 1324.560 ;
    END
  END io_fdi_plConfig_bits[27]
  PIN io_fdi_plConfig_bits[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1.000 264.410 4.000 ;
    END
  END io_fdi_plConfig_bits[28]
  PIN io_fdi_plConfig_bits[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1321.560 364.230 1324.560 ;
    END
  END io_fdi_plConfig_bits[29]
  PIN io_fdi_plConfig_bits[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 822.840 4.000 823.440 ;
    END
  END io_fdi_plConfig_bits[2]
  PIN io_fdi_plConfig_bits[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1190.040 1313.840 1190.640 ;
    END
  END io_fdi_plConfig_bits[30]
  PIN io_fdi_plConfig_bits[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1057.440 1313.840 1058.040 ;
    END
  END io_fdi_plConfig_bits[31]
  PIN io_fdi_plConfig_bits[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 765.040 1313.840 765.640 ;
    END
  END io_fdi_plConfig_bits[3]
  PIN io_fdi_plConfig_bits[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 1.000 821.470 4.000 ;
    END
  END io_fdi_plConfig_bits[4]
  PIN io_fdi_plConfig_bits[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1321.560 663.690 1324.560 ;
    END
  END io_fdi_plConfig_bits[5]
  PIN io_fdi_plConfig_bits[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1.000 19.690 4.000 ;
    END
  END io_fdi_plConfig_bits[6]
  PIN io_fdi_plConfig_bits[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 1.000 357.790 4.000 ;
    END
  END io_fdi_plConfig_bits[7]
  PIN io_fdi_plConfig_bits[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1321.560 119.510 1324.560 ;
    END
  END io_fdi_plConfig_bits[8]
  PIN io_fdi_plConfig_bits[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1321.560 109.850 1324.560 ;
    END
  END io_fdi_plConfig_bits[9]
  PIN io_fdi_plConfig_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1.000 985.690 4.000 ;
    END
  END io_fdi_plConfig_valid
  PIN io_fdi_plData_bits[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 125.840 1313.840 126.440 ;
    END
  END io_fdi_plData_bits[0]
  PIN io_fdi_plData_bits[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 748.040 4.000 748.640 ;
    END
  END io_fdi_plData_bits[10]
  PIN io_fdi_plData_bits[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1.000 1178.890 4.000 ;
    END
  END io_fdi_plData_bits[11]
  PIN io_fdi_plData_bits[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 918.040 1313.840 918.640 ;
    END
  END io_fdi_plData_bits[12]
  PIN io_fdi_plData_bits[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 1.000 872.990 4.000 ;
    END
  END io_fdi_plData_bits[13]
  PIN io_fdi_plData_bits[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1321.560 293.390 1324.560 ;
    END
  END io_fdi_plData_bits[14]
  PIN io_fdi_plData_bits[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1321.560 335.250 1324.560 ;
    END
  END io_fdi_plData_bits[15]
  PIN io_fdi_plData_bits[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1016.640 4.000 1017.240 ;
    END
  END io_fdi_plData_bits[16]
  PIN io_fdi_plData_bits[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 91.840 1313.840 92.440 ;
    END
  END io_fdi_plData_bits[17]
  PIN io_fdi_plData_bits[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 10.240 4.000 10.840 ;
    END
  END io_fdi_plData_bits[18]
  PIN io_fdi_plData_bits[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 853.440 4.000 854.040 ;
    END
  END io_fdi_plData_bits[19]
  PIN io_fdi_plData_bits[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 74.840 4.000 75.440 ;
    END
  END io_fdi_plData_bits[1]
  PIN io_fdi_plData_bits[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1159.440 4.000 1160.040 ;
    END
  END io_fdi_plData_bits[20]
  PIN io_fdi_plData_bits[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 656.240 1313.840 656.840 ;
    END
  END io_fdi_plData_bits[21]
  PIN io_fdi_plData_bits[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 1321.560 406.090 1324.560 ;
    END
  END io_fdi_plData_bits[22]
  PIN io_fdi_plData_bits[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 1.000 1159.570 4.000 ;
    END
  END io_fdi_plData_bits[23]
  PIN io_fdi_plData_bits[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 829.640 1313.840 830.240 ;
    END
  END io_fdi_plData_bits[24]
  PIN io_fdi_plData_bits[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1.000 676.570 4.000 ;
    END
  END io_fdi_plData_bits[25]
  PIN io_fdi_plData_bits[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 190.440 1313.840 191.040 ;
    END
  END io_fdi_plData_bits[26]
  PIN io_fdi_plData_bits[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1321.560 776.390 1324.560 ;
    END
  END io_fdi_plData_bits[27]
  PIN io_fdi_plData_bits[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1203.640 4.000 1204.240 ;
    END
  END io_fdi_plData_bits[28]
  PIN io_fdi_plData_bits[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1.000 441.510 4.000 ;
    END
  END io_fdi_plData_bits[29]
  PIN io_fdi_plData_bits[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1.000 695.890 4.000 ;
    END
  END io_fdi_plData_bits[2]
  PIN io_fdi_plData_bits[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1321.560 200.010 1324.560 ;
    END
  END io_fdi_plData_bits[30]
  PIN io_fdi_plData_bits[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1.000 151.710 4.000 ;
    END
  END io_fdi_plData_bits[31]
  PIN io_fdi_plData_bits[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 1321.560 541.330 1324.560 ;
    END
  END io_fdi_plData_bits[32]
  PIN io_fdi_plData_bits[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 1.000 1149.910 4.000 ;
    END
  END io_fdi_plData_bits[33]
  PIN io_fdi_plData_bits[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 1.000 470.490 4.000 ;
    END
  END io_fdi_plData_bits[34]
  PIN io_fdi_plData_bits[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 724.240 4.000 724.840 ;
    END
  END io_fdi_plData_bits[35]
  PIN io_fdi_plData_bits[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 1321.560 827.910 1324.560 ;
    END
  END io_fdi_plData_bits[36]
  PIN io_fdi_plData_bits[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 333.240 4.000 333.840 ;
    END
  END io_fdi_plData_bits[37]
  PIN io_fdi_plData_bits[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 1.000 976.030 4.000 ;
    END
  END io_fdi_plData_bits[38]
  PIN io_fdi_plData_bits[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 530.440 4.000 531.040 ;
    END
  END io_fdi_plData_bits[39]
  PIN io_fdi_plData_bits[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 1321.560 1175.670 1324.560 ;
    END
  END io_fdi_plData_bits[3]
  PIN io_fdi_plData_bits[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 421.640 4.000 422.240 ;
    END
  END io_fdi_plData_bits[40]
  PIN io_fdi_plData_bits[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1.000 480.150 4.000 ;
    END
  END io_fdi_plData_bits[41]
  PIN io_fdi_plData_bits[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 1.000 1291.590 4.000 ;
    END
  END io_fdi_plData_bits[42]
  PIN io_fdi_plData_bits[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 581.440 1313.840 582.040 ;
    END
  END io_fdi_plData_bits[43]
  PIN io_fdi_plData_bits[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 1321.560 1291.590 1324.560 ;
    END
  END io_fdi_plData_bits[44]
  PIN io_fdi_plData_bits[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 873.840 1313.840 874.440 ;
    END
  END io_fdi_plData_bits[45]
  PIN io_fdi_plData_bits[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 802.440 4.000 803.040 ;
    END
  END io_fdi_plData_bits[46]
  PIN io_fdi_plData_bits[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 411.440 4.000 412.040 ;
    END
  END io_fdi_plData_bits[47]
  PIN io_fdi_plData_bits[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 1321.560 1207.870 1324.560 ;
    END
  END io_fdi_plData_bits[48]
  PIN io_fdi_plData_bits[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1135.640 4.000 1136.240 ;
    END
  END io_fdi_plData_bits[49]
  PIN io_fdi_plData_bits[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1298.840 1313.840 1299.440 ;
    END
  END io_fdi_plData_bits[4]
  PIN io_fdi_plData_bits[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1321.560 621.830 1324.560 ;
    END
  END io_fdi_plData_bits[50]
  PIN io_fdi_plData_bits[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1234.240 4.000 1234.840 ;
    END
  END io_fdi_plData_bits[51]
  PIN io_fdi_plData_bits[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1321.560 766.730 1324.560 ;
    END
  END io_fdi_plData_bits[52]
  PIN io_fdi_plData_bits[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1321.560 415.750 1324.560 ;
    END
  END io_fdi_plData_bits[53]
  PIN io_fdi_plData_bits[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1321.560 795.710 1324.560 ;
    END
  END io_fdi_plData_bits[54]
  PIN io_fdi_plData_bits[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 1321.560 1227.190 1324.560 ;
    END
  END io_fdi_plData_bits[55]
  PIN io_fdi_plData_bits[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 465.840 4.000 466.440 ;
    END
  END io_fdi_plData_bits[56]
  PIN io_fdi_plData_bits[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1321.560 612.170 1324.560 ;
    END
  END io_fdi_plData_bits[57]
  PIN io_fdi_plData_bits[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1321.560 283.730 1324.560 ;
    END
  END io_fdi_plData_bits[58]
  PIN io_fdi_plData_bits[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1321.560 428.630 1324.560 ;
    END
  END io_fdi_plData_bits[59]
  PIN io_fdi_plData_bits[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1.000 563.870 4.000 ;
    END
  END io_fdi_plData_bits[5]
  PIN io_fdi_plData_bits[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 1.000 554.210 4.000 ;
    END
  END io_fdi_plData_bits[60]
  PIN io_fdi_plData_bits[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1275.040 1313.840 1275.640 ;
    END
  END io_fdi_plData_bits[61]
  PIN io_fdi_plData_bits[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1.000 573.530 4.000 ;
    END
  END io_fdi_plData_bits[62]
  PIN io_fdi_plData_bits[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 669.840 4.000 670.440 ;
    END
  END io_fdi_plData_bits[63]
  PIN io_fdi_plData_bits[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 921.440 4.000 922.040 ;
    END
  END io_fdi_plData_bits[6]
  PIN io_fdi_plData_bits[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 887.440 4.000 888.040 ;
    END
  END io_fdi_plData_bits[7]
  PIN io_fdi_plData_bits[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 1321.560 303.050 1324.560 ;
    END
  END io_fdi_plData_bits[8]
  PIN io_fdi_plData_bits[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 333.240 1313.840 333.840 ;
    END
  END io_fdi_plData_bits[9]
  PIN io_fdi_plData_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1213.840 4.000 1214.440 ;
    END
  END io_fdi_plData_valid
  PIN io_fdi_plDllpOfc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1321.560 560.650 1324.560 ;
    END
  END io_fdi_plDllpOfc
  PIN io_fdi_plDllp_bits[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 1.000 512.350 4.000 ;
    END
  END io_fdi_plDllp_bits[0]
  PIN io_fdi_plDllp_bits[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 377.440 4.000 378.040 ;
    END
  END io_fdi_plDllp_bits[1]
  PIN io_fdi_plDllp_bits[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 1321.560 377.110 1324.560 ;
    END
  END io_fdi_plDllp_bits[2]
  PIN io_fdi_plDllp_bits[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 1321.560 509.130 1324.560 ;
    END
  END io_fdi_plDllp_bits[3]
  PIN io_fdi_plDllp_bits[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 1321.560 1301.250 1324.560 ;
    END
  END io_fdi_plDllp_bits[4]
  PIN io_fdi_plDllp_bits[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1321.560 695.890 1324.560 ;
    END
  END io_fdi_plDllp_bits[5]
  PIN io_fdi_plDllp_bits[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 1.000 644.370 4.000 ;
    END
  END io_fdi_plDllp_bits[6]
  PIN io_fdi_plDllp_bits[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 1321.560 1278.710 1324.560 ;
    END
  END io_fdi_plDllp_bits[7]
  PIN io_fdi_plDllp_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 387.640 1313.840 388.240 ;
    END
  END io_fdi_plDllp_valid
  PIN io_fdi_plError
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1.000 544.550 4.000 ;
    END
  END io_fdi_plError
  PIN io_fdi_plFlitCancel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 1.000 1188.550 4.000 ;
    END
  END io_fdi_plFlitCancel
  PIN io_fdi_plInbandPres
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 30.640 4.000 31.240 ;
    END
  END io_fdi_plInbandPres
  PIN io_fdi_plLinkWidth[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 6.840 1313.840 7.440 ;
    END
  END io_fdi_plLinkWidth[0]
  PIN io_fdi_plLinkWidth[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1288.640 4.000 1289.240 ;
    END
  END io_fdi_plLinkWidth[1]
  PIN io_fdi_plLinkWidth[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.640 4.000 184.240 ;
    END
  END io_fdi_plLinkWidth[2]
  PIN io_fdi_plNfError
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 1321.560 232.210 1324.560 ;
    END
  END io_fdi_plNfError
  PIN io_fdi_plPhyInL1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 214.240 4.000 214.840 ;
    END
  END io_fdi_plPhyInL1
  PIN io_fdi_plPhyInL2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 907.840 1313.840 908.440 ;
    END
  END io_fdi_plPhyInL2
  PIN io_fdi_plPhyInRecenter
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 1.000 892.310 4.000 ;
    END
  END io_fdi_plPhyInRecenter
  PIN io_fdi_plProtocolFlitFormat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 809.240 1313.840 809.840 ;
    END
  END io_fdi_plProtocolFlitFormat[0]
  PIN io_fdi_plProtocolFlitFormat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 302.640 4.000 303.240 ;
    END
  END io_fdi_plProtocolFlitFormat[1]
  PIN io_fdi_plProtocolFlitFormat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1321.560 499.470 1324.560 ;
    END
  END io_fdi_plProtocolFlitFormat[2]
  PIN io_fdi_plProtocolValid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 374.040 1313.840 374.640 ;
    END
  END io_fdi_plProtocolValid
  PIN io_fdi_plProtocol[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1.000 583.190 4.000 ;
    END
  END io_fdi_plProtocol[0]
  PIN io_fdi_plProtocol[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 193.840 4.000 194.440 ;
    END
  END io_fdi_plProtocol[1]
  PIN io_fdi_plProtocol[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1321.560 1104.830 1324.560 ;
    END
  END io_fdi_plProtocol[2]
  PIN io_fdi_plRetimerCrd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1321.560 1240.070 1324.560 ;
    END
  END io_fdi_plRetimerCrd
  PIN io_fdi_plRxActiveReq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 1321.560 1085.510 1324.560 ;
    END
  END io_fdi_plRxActiveReq
  PIN io_fdi_plSpeedMode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 40.840 4.000 41.440 ;
    END
  END io_fdi_plSpeedMode[0]
  PIN io_fdi_plSpeedMode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1122.040 1313.840 1122.640 ;
    END
  END io_fdi_plSpeedMode[1]
  PIN io_fdi_plSpeedMode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1.000 315.930 4.000 ;
    END
  END io_fdi_plSpeedMode[2]
  PIN io_fdi_plStallReq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1321.560 325.590 1324.560 ;
    END
  END io_fdi_plStallReq
  PIN io_fdi_plStateStatus[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1040.440 4.000 1041.040 ;
    END
  END io_fdi_plStateStatus[0]
  PIN io_fdi_plStateStatus[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 1321.560 837.570 1324.560 ;
    END
  END io_fdi_plStateStatus[1]
  PIN io_fdi_plStateStatus[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1135.640 1313.840 1136.240 ;
    END
  END io_fdi_plStateStatus[2]
  PIN io_fdi_plStateStatus[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 1321.560 1114.490 1324.560 ;
    END
  END io_fdi_plStateStatus[3]
  PIN io_fdi_plStream_protoStack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1.000 1127.370 4.000 ;
    END
  END io_fdi_plStream_protoStack
  PIN io_fdi_plStream_protoType[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1.000 502.690 4.000 ;
    END
  END io_fdi_plStream_protoType[0]
  PIN io_fdi_plStream_protoType[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1190.040 4.000 1190.640 ;
    END
  END io_fdi_plStream_protoType[1]
  PIN io_fdi_plStream_protoType[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 367.240 4.000 367.840 ;
    END
  END io_fdi_plStream_protoType[2]
  PIN io_fdi_plTrainError
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 1321.560 592.850 1324.560 ;
    END
  END io_fdi_plTrainError
  PIN io_fdi_plWakeAck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1166.240 1313.840 1166.840 ;
    END
  END io_fdi_plWakeAck
  PIN io_rdi_lpClkAck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 703.840 4.000 704.440 ;
    END
  END io_rdi_lpClkAck
  PIN io_rdi_lpConfigCredit
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1321.560 1062.970 1324.560 ;
    END
  END io_rdi_lpConfigCredit
  PIN io_rdi_lpConfig_bits[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 1321.560 1011.450 1324.560 ;
    END
  END io_rdi_lpConfig_bits[0]
  PIN io_rdi_lpConfig_bits[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1321.560 489.810 1324.560 ;
    END
  END io_rdi_lpConfig_bits[10]
  PIN io_rdi_lpConfig_bits[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 472.640 1313.840 473.240 ;
    END
  END io_rdi_lpConfig_bits[11]
  PIN io_rdi_lpConfig_bits[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1321.560 1249.730 1324.560 ;
    END
  END io_rdi_lpConfig_bits[12]
  PIN io_rdi_lpConfig_bits[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1254.640 1313.840 1255.240 ;
    END
  END io_rdi_lpConfig_bits[13]
  PIN io_rdi_lpConfig_bits[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1.000 451.170 4.000 ;
    END
  END io_rdi_lpConfig_bits[14]
  PIN io_rdi_lpConfig_bits[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 710.640 1313.840 711.240 ;
    END
  END io_rdi_lpConfig_bits[15]
  PIN io_rdi_lpConfig_bits[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 1.000 831.130 4.000 ;
    END
  END io_rdi_lpConfig_bits[16]
  PIN io_rdi_lpConfig_bits[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 428.440 1313.840 429.040 ;
    END
  END io_rdi_lpConfig_bits[17]
  PIN io_rdi_lpConfig_bits[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 1321.560 457.610 1324.560 ;
    END
  END io_rdi_lpConfig_bits[18]
  PIN io_rdi_lpConfig_bits[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 659.640 4.000 660.240 ;
    END
  END io_rdi_lpConfig_bits[19]
  PIN io_rdi_lpConfig_bits[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1.000 666.910 4.000 ;
    END
  END io_rdi_lpConfig_bits[1]
  PIN io_rdi_lpConfig_bits[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 1.000 592.850 4.000 ;
    END
  END io_rdi_lpConfig_bits[20]
  PIN io_rdi_lpConfig_bits[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 948.640 1313.840 949.240 ;
    END
  END io_rdi_lpConfig_bits[21]
  PIN io_rdi_lpConfig_bits[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 289.040 1313.840 289.640 ;
    END
  END io_rdi_lpConfig_bits[22]
  PIN io_rdi_lpConfig_bits[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 1.000 1211.090 4.000 ;
    END
  END io_rdi_lpConfig_bits[23]
  PIN io_rdi_lpConfig_bits[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 506.640 1313.840 507.240 ;
    END
  END io_rdi_lpConfig_bits[24]
  PIN io_rdi_lpConfig_bits[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 931.640 4.000 932.240 ;
    END
  END io_rdi_lpConfig_bits[25]
  PIN io_rdi_lpConfig_bits[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 540.640 4.000 541.240 ;
    END
  END io_rdi_lpConfig_bits[26]
  PIN io_rdi_lpConfig_bits[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 1321.560 1166.010 1324.560 ;
    END
  END io_rdi_lpConfig_bits[27]
  PIN io_rdi_lpConfig_bits[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 941.840 4.000 942.440 ;
    END
  END io_rdi_lpConfig_bits[28]
  PIN io_rdi_lpConfig_bits[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 234.640 1313.840 235.240 ;
    END
  END io_rdi_lpConfig_bits[29]
  PIN io_rdi_lpConfig_bits[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 506.640 4.000 507.240 ;
    END
  END io_rdi_lpConfig_bits[2]
  PIN io_rdi_lpConfig_bits[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1.000 953.490 4.000 ;
    END
  END io_rdi_lpConfig_bits[30]
  PIN io_rdi_lpConfig_bits[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 136.040 1313.840 136.640 ;
    END
  END io_rdi_lpConfig_bits[31]
  PIN io_rdi_lpConfig_bits[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 669.840 1313.840 670.440 ;
    END
  END io_rdi_lpConfig_bits[3]
  PIN io_rdi_lpConfig_bits[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1321.560 1137.030 1324.560 ;
    END
  END io_rdi_lpConfig_bits[4]
  PIN io_rdi_lpConfig_bits[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 224.440 4.000 225.040 ;
    END
  END io_rdi_lpConfig_bits[5]
  PIN io_rdi_lpConfig_bits[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1169.640 4.000 1170.240 ;
    END
  END io_rdi_lpConfig_bits[6]
  PIN io_rdi_lpConfig_bits[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1321.560 447.950 1324.560 ;
    END
  END io_rdi_lpConfig_bits[7]
  PIN io_rdi_lpConfig_bits[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1321.560 48.670 1324.560 ;
    END
  END io_rdi_lpConfig_bits[8]
  PIN io_rdi_lpConfig_bits[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1.000 71.210 4.000 ;
    END
  END io_rdi_lpConfig_bits[9]
  PIN io_rdi_lpConfig_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 1.000 338.470 4.000 ;
    END
  END io_rdi_lpConfig_valid
  PIN io_rdi_lpData_bits[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 27.240 1313.840 27.840 ;
    END
  END io_rdi_lpData_bits[0]
  PIN io_rdi_lpData_bits[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 972.440 1313.840 973.040 ;
    END
  END io_rdi_lpData_bits[10]
  PIN io_rdi_lpData_bits[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 952.040 4.000 952.640 ;
    END
  END io_rdi_lpData_bits[11]
  PIN io_rdi_lpData_bits[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1081.240 4.000 1081.840 ;
    END
  END io_rdi_lpData_bits[12]
  PIN io_rdi_lpData_bits[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1321.560 58.330 1324.560 ;
    END
  END io_rdi_lpData_bits[13]
  PIN io_rdi_lpData_bits[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1.000 808.590 4.000 ;
    END
  END io_rdi_lpData_bits[14]
  PIN io_rdi_lpData_bits[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 1321.560 644.370 1324.560 ;
    END
  END io_rdi_lpData_bits[15]
  PIN io_rdi_lpData_bits[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1071.040 4.000 1071.640 ;
    END
  END io_rdi_lpData_bits[16]
  PIN io_rdi_lpData_bits[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 516.840 1313.840 517.440 ;
    END
  END io_rdi_lpData_bits[17]
  PIN io_rdi_lpData_bits[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1081.240 1313.840 1081.840 ;
    END
  END io_rdi_lpData_bits[18]
  PIN io_rdi_lpData_bits[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1220.640 1313.840 1221.240 ;
    END
  END io_rdi_lpData_bits[19]
  PIN io_rdi_lpData_bits[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 907.840 4.000 908.440 ;
    END
  END io_rdi_lpData_bits[1]
  PIN io_rdi_lpData_bits[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1071.040 1313.840 1071.640 ;
    END
  END io_rdi_lpData_bits[20]
  PIN io_rdi_lpData_bits[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1321.560 705.550 1324.560 ;
    END
  END io_rdi_lpData_bits[21]
  PIN io_rdi_lpData_bits[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 1.000 389.990 4.000 ;
    END
  END io_rdi_lpData_bits[22]
  PIN io_rdi_lpData_bits[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1321.560 467.270 1324.560 ;
    END
  END io_rdi_lpData_bits[23]
  PIN io_rdi_lpData_bits[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 255.040 1313.840 255.640 ;
    END
  END io_rdi_lpData_bits[24]
  PIN io_rdi_lpData_bits[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 571.240 1313.840 571.840 ;
    END
  END io_rdi_lpData_bits[25]
  PIN io_rdi_lpData_bits[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 159.840 4.000 160.440 ;
    END
  END io_rdi_lpData_bits[26]
  PIN io_rdi_lpData_bits[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 574.640 4.000 575.240 ;
    END
  END io_rdi_lpData_bits[27]
  PIN io_rdi_lpData_bits[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 863.640 1313.840 864.240 ;
    END
  END io_rdi_lpData_bits[28]
  PIN io_rdi_lpData_bits[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 700.440 1313.840 701.040 ;
    END
  END io_rdi_lpData_bits[29]
  PIN io_rdi_lpData_bits[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1210.440 1313.840 1211.040 ;
    END
  END io_rdi_lpData_bits[2]
  PIN io_rdi_lpData_bits[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 105.440 4.000 106.040 ;
    END
  END io_rdi_lpData_bits[30]
  PIN io_rdi_lpData_bits[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1.000 1098.390 4.000 ;
    END
  END io_rdi_lpData_bits[31]
  PIN io_rdi_lpData_bits[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1016.640 1313.840 1017.240 ;
    END
  END io_rdi_lpData_bits[32]
  PIN io_rdi_lpData_bits[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1.000 1056.530 4.000 ;
    END
  END io_rdi_lpData_bits[33]
  PIN io_rdi_lpData_bits[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1321.560 354.570 1324.560 ;
    END
  END io_rdi_lpData_bits[34]
  PIN io_rdi_lpData_bits[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 476.040 4.000 476.640 ;
    END
  END io_rdi_lpData_bits[35]
  PIN io_rdi_lpData_bits[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 1.000 328.810 4.000 ;
    END
  END io_rdi_lpData_bits[36]
  PIN io_rdi_lpData_bits[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 1.000 1140.250 4.000 ;
    END
  END io_rdi_lpData_bits[37]
  PIN io_rdi_lpData_bits[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 244.840 1313.840 245.440 ;
    END
  END io_rdi_lpData_bits[38]
  PIN io_rdi_lpData_bits[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1030.240 4.000 1030.840 ;
    END
  END io_rdi_lpData_bits[39]
  PIN io_rdi_lpData_bits[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 550.840 4.000 551.440 ;
    END
  END io_rdi_lpData_bits[3]
  PIN io_rdi_lpData_bits[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1321.560 129.170 1324.560 ;
    END
  END io_rdi_lpData_bits[40]
  PIN io_rdi_lpData_bits[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1321.560 26.130 1324.560 ;
    END
  END io_rdi_lpData_bits[41]
  PIN io_rdi_lpData_bits[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1.000 399.650 4.000 ;
    END
  END io_rdi_lpData_bits[42]
  PIN io_rdi_lpData_bits[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1026.840 1313.840 1027.440 ;
    END
  END io_rdi_lpData_bits[43]
  PIN io_rdi_lpData_bits[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 1.000 1262.610 4.000 ;
    END
  END io_rdi_lpData_bits[44]
  PIN io_rdi_lpData_bits[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 1321.560 602.510 1324.560 ;
    END
  END io_rdi_lpData_bits[45]
  PIN io_rdi_lpData_bits[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 1.000 254.750 4.000 ;
    END
  END io_rdi_lpData_bits[46]
  PIN io_rdi_lpData_bits[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 884.040 1313.840 884.640 ;
    END
  END io_rdi_lpData_bits[47]
  PIN io_rdi_lpData_bits[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1321.560 1124.150 1324.560 ;
    END
  END io_rdi_lpData_bits[48]
  PIN io_rdi_lpData_bits[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1321.560 1053.310 1324.560 ;
    END
  END io_rdi_lpData_bits[49]
  PIN io_rdi_lpData_bits[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 1321.560 1269.050 1324.560 ;
    END
  END io_rdi_lpData_bits[4]
  PIN io_rdi_lpData_bits[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1319.240 1313.840 1319.840 ;
    END
  END io_rdi_lpData_bits[50]
  PIN io_rdi_lpData_bits[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1309.040 1313.840 1309.640 ;
    END
  END io_rdi_lpData_bits[51]
  PIN io_rdi_lpData_bits[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1.000 718.430 4.000 ;
    END
  END io_rdi_lpData_bits[52]
  PIN io_rdi_lpData_bits[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 1321.560 921.290 1324.560 ;
    END
  END io_rdi_lpData_bits[53]
  PIN io_rdi_lpData_bits[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 51.040 4.000 51.640 ;
    END
  END io_rdi_lpData_bits[54]
  PIN io_rdi_lpData_bits[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1.000 10.030 4.000 ;
    END
  END io_rdi_lpData_bits[55]
  PIN io_rdi_lpData_bits[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 520.240 4.000 520.840 ;
    END
  END io_rdi_lpData_bits[56]
  PIN io_rdi_lpData_bits[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1.000 728.090 4.000 ;
    END
  END io_rdi_lpData_bits[57]
  PIN io_rdi_lpData_bits[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 323.040 4.000 323.640 ;
    END
  END io_rdi_lpData_bits[58]
  PIN io_rdi_lpData_bits[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 561.040 4.000 561.640 ;
    END
  END io_rdi_lpData_bits[59]
  PIN io_rdi_lpData_bits[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 268.640 1313.840 269.240 ;
    END
  END io_rdi_lpData_bits[5]
  PIN io_rdi_lpData_bits[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1321.560 212.890 1324.560 ;
    END
  END io_rdi_lpData_bits[60]
  PIN io_rdi_lpData_bits[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 714.040 4.000 714.640 ;
    END
  END io_rdi_lpData_bits[61]
  PIN io_rdi_lpData_bits[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 238.040 4.000 238.640 ;
    END
  END io_rdi_lpData_bits[62]
  PIN io_rdi_lpData_bits[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1.000 615.390 4.000 ;
    END
  END io_rdi_lpData_bits[63]
  PIN io_rdi_lpData_bits[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 85.040 4.000 85.640 ;
    END
  END io_rdi_lpData_bits[6]
  PIN io_rdi_lpData_bits[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 1.000 1117.710 4.000 ;
    END
  END io_rdi_lpData_bits[7]
  PIN io_rdi_lpData_bits[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1.000 531.670 4.000 ;
    END
  END io_rdi_lpData_bits[8]
  PIN io_rdi_lpData_bits[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1321.560 6.810 1324.560 ;
    END
  END io_rdi_lpData_bits[9]
  PIN io_rdi_lpData_irdy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1254.640 4.000 1255.240 ;
    END
  END io_rdi_lpData_irdy
  PIN io_rdi_lpData_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1047.240 1313.840 1047.840 ;
    END
  END io_rdi_lpData_ready
  PIN io_rdi_lpData_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 1.000 1066.190 4.000 ;
    END
  END io_rdi_lpData_valid
  PIN io_rdi_lpLinkError
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1321.560 180.690 1324.560 ;
    END
  END io_rdi_lpLinkError
  PIN io_rdi_lpRetimerCrd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 486.240 4.000 486.840 ;
    END
  END io_rdi_lpRetimerCrd
  PIN io_rdi_lpStallAck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 992.840 1313.840 993.440 ;
    END
  END io_rdi_lpStallAck
  PIN io_rdi_lpStateReq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1321.560 683.010 1324.560 ;
    END
  END io_rdi_lpStateReq[0]
  PIN io_rdi_lpStateReq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 819.440 1313.840 820.040 ;
    END
  END io_rdi_lpStateReq[1]
  PIN io_rdi_lpStateReq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 843.240 4.000 843.840 ;
    END
  END io_rdi_lpStateReq[2]
  PIN io_rdi_lpStateReq[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1321.560 982.470 1324.560 ;
    END
  END io_rdi_lpStateReq[3]
  PIN io_rdi_lpWakeReq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 214.240 1313.840 214.840 ;
    END
  END io_rdi_lpWakeReq
  PIN io_rdi_plClkReq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1321.560 579.970 1324.560 ;
    END
  END io_rdi_plClkReq
  PIN io_rdi_plConfigCredit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 1.000 1272.270 4.000 ;
    END
  END io_rdi_plConfigCredit
  PIN io_rdi_plConfig_bits[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1321.560 100.190 1324.560 ;
    END
  END io_rdi_plConfig_bits[0]
  PIN io_rdi_plConfig_bits[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1.000 174.250 4.000 ;
    END
  END io_rdi_plConfig_bits[10]
  PIN io_rdi_plConfig_bits[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 788.840 1313.840 789.440 ;
    END
  END io_rdi_plConfig_bits[11]
  PIN io_rdi_plConfig_bits[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 975.840 4.000 976.440 ;
    END
  END io_rdi_plConfig_bits[12]
  PIN io_rdi_plConfig_bits[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1050.640 4.000 1051.240 ;
    END
  END io_rdi_plConfig_bits[13]
  PIN io_rdi_plConfig_bits[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1.000 348.130 4.000 ;
    END
  END io_rdi_plConfig_bits[14]
  PIN io_rdi_plConfig_bits[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 734.440 4.000 735.040 ;
    END
  END io_rdi_plConfig_bits[15]
  PIN io_rdi_plConfig_bits[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1321.560 190.350 1324.560 ;
    END
  END io_rdi_plConfig_bits[16]
  PIN io_rdi_plConfig_bits[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1321.560 959.930 1324.560 ;
    END
  END io_rdi_plConfig_bits[17]
  PIN io_rdi_plConfig_bits[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1145.840 1313.840 1146.440 ;
    END
  END io_rdi_plConfig_bits[18]
  PIN io_rdi_plConfig_bits[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1321.560 138.830 1324.560 ;
    END
  END io_rdi_plConfig_bits[19]
  PIN io_rdi_plConfig_bits[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1321.560 264.410 1324.560 ;
    END
  END io_rdi_plConfig_bits[1]
  PIN io_rdi_plConfig_bits[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 299.240 1313.840 299.840 ;
    END
  END io_rdi_plConfig_bits[20]
  PIN io_rdi_plConfig_bits[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1321.560 67.990 1324.560 ;
    END
  END io_rdi_plConfig_bits[21]
  PIN io_rdi_plConfig_bits[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 547.440 1313.840 548.040 ;
    END
  END io_rdi_plConfig_bits[22]
  PIN io_rdi_plConfig_bits[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 996.240 4.000 996.840 ;
    END
  END io_rdi_plConfig_bits[23]
  PIN io_rdi_plConfig_bits[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 1321.560 438.290 1324.560 ;
    END
  END io_rdi_plConfig_bits[24]
  PIN io_rdi_plConfig_bits[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1224.040 4.000 1224.640 ;
    END
  END io_rdi_plConfig_bits[25]
  PIN io_rdi_plConfig_bits[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1.000 122.730 4.000 ;
    END
  END io_rdi_plConfig_bits[26]
  PIN io_rdi_plConfig_bits[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 605.240 4.000 605.840 ;
    END
  END io_rdi_plConfig_bits[27]
  PIN io_rdi_plConfig_bits[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 278.840 4.000 279.440 ;
    END
  END io_rdi_plConfig_bits[28]
  PIN io_rdi_plConfig_bits[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1003.040 1313.840 1003.640 ;
    END
  END io_rdi_plConfig_bits[29]
  PIN io_rdi_plConfig_bits[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1.000 860.110 4.000 ;
    END
  END io_rdi_plConfig_bits[2]
  PIN io_rdi_plConfig_bits[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 897.640 1313.840 898.240 ;
    END
  END io_rdi_plConfig_bits[30]
  PIN io_rdi_plConfig_bits[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 482.840 1313.840 483.440 ;
    END
  END io_rdi_plConfig_bits[31]
  PIN io_rdi_plConfig_bits[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 1.000 1304.470 4.000 ;
    END
  END io_rdi_plConfig_bits[3]
  PIN io_rdi_plConfig_bits[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1321.560 715.210 1324.560 ;
    END
  END io_rdi_plConfig_bits[4]
  PIN io_rdi_plConfig_bits[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1321.560 1095.170 1324.560 ;
    END
  END io_rdi_plConfig_bits[5]
  PIN io_rdi_plConfig_bits[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 1.000 769.950 4.000 ;
    END
  END io_rdi_plConfig_bits[6]
  PIN io_rdi_plConfig_bits[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1.000 1088.730 4.000 ;
    END
  END io_rdi_plConfig_bits[7]
  PIN io_rdi_plConfig_bits[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 353.640 1313.840 354.240 ;
    END
  END io_rdi_plConfig_bits[8]
  PIN io_rdi_plConfig_bits[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1321.560 16.470 1324.560 ;
    END
  END io_rdi_plConfig_bits[9]
  PIN io_rdi_plConfig_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1.000 737.750 4.000 ;
    END
  END io_rdi_plConfig_valid
  PIN io_rdi_plCorrectableError
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 1.000 142.050 4.000 ;
    END
  END io_rdi_plCorrectableError
  PIN io_rdi_plData_bits[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 768.440 4.000 769.040 ;
    END
  END io_rdi_plData_bits[0]
  PIN io_rdi_plData_bits[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 625.640 4.000 626.240 ;
    END
  END io_rdi_plData_bits[10]
  PIN io_rdi_plData_bits[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 1321.560 1259.390 1324.560 ;
    END
  END io_rdi_plData_bits[11]
  PIN io_rdi_plData_bits[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 1.000 522.010 4.000 ;
    END
  END io_rdi_plData_bits[12]
  PIN io_rdi_plData_bits[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 1321.560 930.950 1324.560 ;
    END
  END io_rdi_plData_bits[13]
  PIN io_rdi_plData_bits[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 625.640 1313.840 626.240 ;
    END
  END io_rdi_plData_bits[14]
  PIN io_rdi_plData_bits[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1.000 1046.870 4.000 ;
    END
  END io_rdi_plData_bits[15]
  PIN io_rdi_plData_bits[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 346.840 4.000 347.440 ;
    END
  END io_rdi_plData_bits[16]
  PIN io_rdi_plData_bits[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 1.000 1005.010 4.000 ;
    END
  END io_rdi_plData_bits[17]
  PIN io_rdi_plData_bits[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1.000 418.970 4.000 ;
    END
  END io_rdi_plData_bits[18]
  PIN io_rdi_plData_bits[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1.000 61.550 4.000 ;
    END
  END io_rdi_plData_bits[19]
  PIN io_rdi_plData_bits[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 17.040 1313.840 17.640 ;
    END
  END io_rdi_plData_bits[1]
  PIN io_rdi_plData_bits[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 397.840 1313.840 398.440 ;
    END
  END io_rdi_plData_bits[20]
  PIN io_rdi_plData_bits[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1321.560 315.930 1324.560 ;
    END
  END io_rdi_plData_bits[21]
  PIN io_rdi_plData_bits[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1244.440 1313.840 1245.040 ;
    END
  END io_rdi_plData_bits[22]
  PIN io_rdi_plData_bits[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 897.640 4.000 898.240 ;
    END
  END io_rdi_plData_bits[23]
  PIN io_rdi_plData_bits[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1006.440 4.000 1007.040 ;
    END
  END io_rdi_plData_bits[24]
  PIN io_rdi_plData_bits[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 962.240 4.000 962.840 ;
    END
  END io_rdi_plData_bits[25]
  PIN io_rdi_plData_bits[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1.000 48.670 4.000 ;
    END
  END io_rdi_plData_bits[26]
  PIN io_rdi_plData_bits[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 139.440 4.000 140.040 ;
    END
  END io_rdi_plData_bits[27]
  PIN io_rdi_plData_bits[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 744.640 1313.840 745.240 ;
    END
  END io_rdi_plData_bits[28]
  PIN io_rdi_plData_bits[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1.000 760.290 4.000 ;
    END
  END io_rdi_plData_bits[29]
  PIN io_rdi_plData_bits[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1321.560 818.250 1324.560 ;
    END
  END io_rdi_plData_bits[2]
  PIN io_rdi_plData_bits[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 1321.560 1146.690 1324.560 ;
    END
  END io_rdi_plData_bits[30]
  PIN io_rdi_plData_bits[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1309.040 4.000 1309.640 ;
    END
  END io_rdi_plData_bits[31]
  PIN io_rdi_plData_bits[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1.000 203.230 4.000 ;
    END
  END io_rdi_plData_bits[32]
  PIN io_rdi_plData_bits[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 853.440 1313.840 854.040 ;
    END
  END io_rdi_plData_bits[33]
  PIN io_rdi_plData_bits[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 1321.560 1188.550 1324.560 ;
    END
  END io_rdi_plData_bits[34]
  PIN io_rdi_plData_bits[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 680.040 4.000 680.640 ;
    END
  END io_rdi_plData_bits[35]
  PIN io_rdi_plData_bits[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1091.440 1313.840 1092.040 ;
    END
  END io_rdi_plData_bits[36]
  PIN io_rdi_plData_bits[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 462.440 1313.840 463.040 ;
    END
  END io_rdi_plData_bits[37]
  PIN io_rdi_plData_bits[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1.000 911.630 4.000 ;
    END
  END io_rdi_plData_bits[38]
  PIN io_rdi_plData_bits[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1321.560 1033.990 1324.560 ;
    END
  END io_rdi_plData_bits[39]
  PIN io_rdi_plData_bits[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1321.560 251.530 1324.560 ;
    END
  END io_rdi_plData_bits[3]
  PIN io_rdi_plData_bits[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1.000 409.310 4.000 ;
    END
  END io_rdi_plData_bits[40]
  PIN io_rdi_plData_bits[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 843.240 1313.840 843.840 ;
    END
  END io_rdi_plData_bits[41]
  PIN io_rdi_plData_bits[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 1.000 1075.850 4.000 ;
    END
  END io_rdi_plData_bits[42]
  PIN io_rdi_plData_bits[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 408.040 1313.840 408.640 ;
    END
  END io_rdi_plData_bits[43]
  PIN io_rdi_plData_bits[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 615.440 4.000 616.040 ;
    END
  END io_rdi_plData_bits[44]
  PIN io_rdi_plData_bits[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 51.040 1313.840 51.640 ;
    END
  END io_rdi_plData_bits[45]
  PIN io_rdi_plData_bits[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1.000 212.890 4.000 ;
    END
  END io_rdi_plData_bits[46]
  PIN io_rdi_plData_bits[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 1.000 657.250 4.000 ;
    END
  END io_rdi_plData_bits[47]
  PIN io_rdi_plData_bits[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 591.640 1313.840 592.240 ;
    END
  END io_rdi_plData_bits[48]
  PIN io_rdi_plData_bits[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 1321.560 992.130 1324.560 ;
    END
  END io_rdi_plData_bits[49]
  PIN io_rdi_plData_bits[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1230.840 1313.840 1231.440 ;
    END
  END io_rdi_plData_bits[4]
  PIN io_rdi_plData_bits[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 61.240 1313.840 61.840 ;
    END
  END io_rdi_plData_bits[50]
  PIN io_rdi_plData_bits[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1.000 100.190 4.000 ;
    END
  END io_rdi_plData_bits[51]
  PIN io_rdi_plData_bits[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 775.240 1313.840 775.840 ;
    END
  END io_rdi_plData_bits[52]
  PIN io_rdi_plData_bits[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1.000 29.350 4.000 ;
    END
  END io_rdi_plData_bits[53]
  PIN io_rdi_plData_bits[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1264.840 1313.840 1265.440 ;
    END
  END io_rdi_plData_bits[54]
  PIN io_rdi_plData_bits[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 1321.560 950.270 1324.560 ;
    END
  END io_rdi_plData_bits[55]
  PIN io_rdi_plData_bits[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 146.240 1313.840 146.840 ;
    END
  END io_rdi_plData_bits[56]
  PIN io_rdi_plData_bits[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1321.560 911.630 1324.560 ;
    END
  END io_rdi_plData_bits[57]
  PIN io_rdi_plData_bits[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 312.840 4.000 313.440 ;
    END
  END io_rdi_plData_bits[58]
  PIN io_rdi_plData_bits[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 357.040 4.000 357.640 ;
    END
  END io_rdi_plData_bits[59]
  PIN io_rdi_plData_bits[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 1.000 882.650 4.000 ;
    END
  END io_rdi_plData_bits[5]
  PIN io_rdi_plData_bits[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END io_rdi_plData_bits[60]
  PIN io_rdi_plData_bits[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1.000 1024.330 4.000 ;
    END
  END io_rdi_plData_bits[61]
  PIN io_rdi_plData_bits[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 595.040 4.000 595.640 ;
    END
  END io_rdi_plData_bits[62]
  PIN io_rdi_plData_bits[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1125.440 4.000 1126.040 ;
    END
  END io_rdi_plData_bits[63]
  PIN io_rdi_plData_bits[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1321.560 344.910 1324.560 ;
    END
  END io_rdi_plData_bits[6]
  PIN io_rdi_plData_bits[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 401.240 4.000 401.840 ;
    END
  END io_rdi_plData_bits[7]
  PIN io_rdi_plData_bits[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 1.000 277.290 4.000 ;
    END
  END io_rdi_plData_bits[8]
  PIN io_rdi_plData_bits[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1.000 90.530 4.000 ;
    END
  END io_rdi_plData_bits[9]
  PIN io_rdi_plData_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1321.560 673.350 1324.560 ;
    END
  END io_rdi_plData_valid
  PIN io_rdi_plError
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1321.560 386.770 1324.560 ;
    END
  END io_rdi_plError
  PIN io_rdi_plInbandPres
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1.000 708.770 4.000 ;
    END
  END io_rdi_plInbandPres
  PIN io_rdi_plLinkWidth[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 1321.560 898.750 1324.560 ;
    END
  END io_rdi_plLinkWidth[0]
  PIN io_rdi_plLinkWidth[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 363.840 1313.840 364.440 ;
    END
  END io_rdi_plLinkWidth[1]
  PIN io_rdi_plLinkWidth[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 867.040 4.000 867.640 ;
    END
  END io_rdi_plLinkWidth[2]
  PIN io_rdi_plNonFatalError
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 1037.040 1313.840 1037.640 ;
    END
  END io_rdi_plNonFatalError
  PIN io_rdi_plPhyInRecenter
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1.000 286.950 4.000 ;
    END
  END io_rdi_plPhyInRecenter
  PIN io_rdi_plRetimerCrd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1.000 493.030 4.000 ;
    END
  END io_rdi_plRetimerCrd
  PIN io_rdi_plSpeedMode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 95.240 4.000 95.840 ;
    END
  END io_rdi_plSpeedMode[0]
  PIN io_rdi_plSpeedMode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 982.640 1313.840 983.240 ;
    END
  END io_rdi_plSpeedMode[1]
  PIN io_rdi_plSpeedMode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1.000 779.610 4.000 ;
    END
  END io_rdi_plSpeedMode[2]
  PIN io_rdi_plStallReq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1321.560 869.770 1324.560 ;
    END
  END io_rdi_plStallReq
  PIN io_rdi_plStateStatus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1321.560 847.230 1324.560 ;
    END
  END io_rdi_plStateStatus[0]
  PIN io_rdi_plStateStatus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1244.440 4.000 1245.040 ;
    END
  END io_rdi_plStateStatus[1]
  PIN io_rdi_plStateStatus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1321.560 161.370 1324.560 ;
    END
  END io_rdi_plStateStatus[2]
  PIN io_rdi_plStateStatus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 1.000 934.170 4.000 ;
    END
  END io_rdi_plStateStatus[3]
  PIN io_rdi_plTrainError
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 292.440 4.000 293.040 ;
    END
  END io_rdi_plTrainError
  PIN io_rdi_plWakeAck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1115.240 4.000 1115.840 ;
    END
  END io_rdi_plWakeAck
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1310.840 635.840 1313.840 636.440 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1309.160 1313.845 ;
      LAYER met1 ;
        RECT 0.070 2.760 1314.610 1317.460 ;
      LAYER met2 ;
        RECT 0.100 1324.840 1314.580 1325.050 ;
        RECT 0.100 1321.280 6.250 1324.840 ;
        RECT 7.090 1321.280 15.910 1324.840 ;
        RECT 16.750 1321.280 25.570 1324.840 ;
        RECT 26.410 1321.280 35.230 1324.840 ;
        RECT 36.070 1321.280 48.110 1324.840 ;
        RECT 48.950 1321.280 57.770 1324.840 ;
        RECT 58.610 1321.280 67.430 1324.840 ;
        RECT 68.270 1321.280 77.090 1324.840 ;
        RECT 77.930 1321.280 86.750 1324.840 ;
        RECT 87.590 1321.280 99.630 1324.840 ;
        RECT 100.470 1321.280 109.290 1324.840 ;
        RECT 110.130 1321.280 118.950 1324.840 ;
        RECT 119.790 1321.280 128.610 1324.840 ;
        RECT 129.450 1321.280 138.270 1324.840 ;
        RECT 139.110 1321.280 147.930 1324.840 ;
        RECT 148.770 1321.280 160.810 1324.840 ;
        RECT 161.650 1321.280 170.470 1324.840 ;
        RECT 171.310 1321.280 180.130 1324.840 ;
        RECT 180.970 1321.280 189.790 1324.840 ;
        RECT 190.630 1321.280 199.450 1324.840 ;
        RECT 200.290 1321.280 212.330 1324.840 ;
        RECT 213.170 1321.280 221.990 1324.840 ;
        RECT 222.830 1321.280 231.650 1324.840 ;
        RECT 232.490 1321.280 241.310 1324.840 ;
        RECT 242.150 1321.280 250.970 1324.840 ;
        RECT 251.810 1321.280 263.850 1324.840 ;
        RECT 264.690 1321.280 273.510 1324.840 ;
        RECT 274.350 1321.280 283.170 1324.840 ;
        RECT 284.010 1321.280 292.830 1324.840 ;
        RECT 293.670 1321.280 302.490 1324.840 ;
        RECT 303.330 1321.280 315.370 1324.840 ;
        RECT 316.210 1321.280 325.030 1324.840 ;
        RECT 325.870 1321.280 334.690 1324.840 ;
        RECT 335.530 1321.280 344.350 1324.840 ;
        RECT 345.190 1321.280 354.010 1324.840 ;
        RECT 354.850 1321.280 363.670 1324.840 ;
        RECT 364.510 1321.280 376.550 1324.840 ;
        RECT 377.390 1321.280 386.210 1324.840 ;
        RECT 387.050 1321.280 395.870 1324.840 ;
        RECT 396.710 1321.280 405.530 1324.840 ;
        RECT 406.370 1321.280 415.190 1324.840 ;
        RECT 416.030 1321.280 428.070 1324.840 ;
        RECT 428.910 1321.280 437.730 1324.840 ;
        RECT 438.570 1321.280 447.390 1324.840 ;
        RECT 448.230 1321.280 457.050 1324.840 ;
        RECT 457.890 1321.280 466.710 1324.840 ;
        RECT 467.550 1321.280 479.590 1324.840 ;
        RECT 480.430 1321.280 489.250 1324.840 ;
        RECT 490.090 1321.280 498.910 1324.840 ;
        RECT 499.750 1321.280 508.570 1324.840 ;
        RECT 509.410 1321.280 518.230 1324.840 ;
        RECT 519.070 1321.280 527.890 1324.840 ;
        RECT 528.730 1321.280 540.770 1324.840 ;
        RECT 541.610 1321.280 550.430 1324.840 ;
        RECT 551.270 1321.280 560.090 1324.840 ;
        RECT 560.930 1321.280 569.750 1324.840 ;
        RECT 570.590 1321.280 579.410 1324.840 ;
        RECT 580.250 1321.280 592.290 1324.840 ;
        RECT 593.130 1321.280 601.950 1324.840 ;
        RECT 602.790 1321.280 611.610 1324.840 ;
        RECT 612.450 1321.280 621.270 1324.840 ;
        RECT 622.110 1321.280 630.930 1324.840 ;
        RECT 631.770 1321.280 643.810 1324.840 ;
        RECT 644.650 1321.280 653.470 1324.840 ;
        RECT 654.310 1321.280 663.130 1324.840 ;
        RECT 663.970 1321.280 672.790 1324.840 ;
        RECT 673.630 1321.280 682.450 1324.840 ;
        RECT 683.290 1321.280 695.330 1324.840 ;
        RECT 696.170 1321.280 704.990 1324.840 ;
        RECT 705.830 1321.280 714.650 1324.840 ;
        RECT 715.490 1321.280 724.310 1324.840 ;
        RECT 725.150 1321.280 733.970 1324.840 ;
        RECT 734.810 1321.280 743.630 1324.840 ;
        RECT 744.470 1321.280 756.510 1324.840 ;
        RECT 757.350 1321.280 766.170 1324.840 ;
        RECT 767.010 1321.280 775.830 1324.840 ;
        RECT 776.670 1321.280 785.490 1324.840 ;
        RECT 786.330 1321.280 795.150 1324.840 ;
        RECT 795.990 1321.280 808.030 1324.840 ;
        RECT 808.870 1321.280 817.690 1324.840 ;
        RECT 818.530 1321.280 827.350 1324.840 ;
        RECT 828.190 1321.280 837.010 1324.840 ;
        RECT 837.850 1321.280 846.670 1324.840 ;
        RECT 847.510 1321.280 859.550 1324.840 ;
        RECT 860.390 1321.280 869.210 1324.840 ;
        RECT 870.050 1321.280 878.870 1324.840 ;
        RECT 879.710 1321.280 888.530 1324.840 ;
        RECT 889.370 1321.280 898.190 1324.840 ;
        RECT 899.030 1321.280 911.070 1324.840 ;
        RECT 911.910 1321.280 920.730 1324.840 ;
        RECT 921.570 1321.280 930.390 1324.840 ;
        RECT 931.230 1321.280 940.050 1324.840 ;
        RECT 940.890 1321.280 949.710 1324.840 ;
        RECT 950.550 1321.280 959.370 1324.840 ;
        RECT 960.210 1321.280 972.250 1324.840 ;
        RECT 973.090 1321.280 981.910 1324.840 ;
        RECT 982.750 1321.280 991.570 1324.840 ;
        RECT 992.410 1321.280 1001.230 1324.840 ;
        RECT 1002.070 1321.280 1010.890 1324.840 ;
        RECT 1011.730 1321.280 1023.770 1324.840 ;
        RECT 1024.610 1321.280 1033.430 1324.840 ;
        RECT 1034.270 1321.280 1043.090 1324.840 ;
        RECT 1043.930 1321.280 1052.750 1324.840 ;
        RECT 1053.590 1321.280 1062.410 1324.840 ;
        RECT 1063.250 1321.280 1075.290 1324.840 ;
        RECT 1076.130 1321.280 1084.950 1324.840 ;
        RECT 1085.790 1321.280 1094.610 1324.840 ;
        RECT 1095.450 1321.280 1104.270 1324.840 ;
        RECT 1105.110 1321.280 1113.930 1324.840 ;
        RECT 1114.770 1321.280 1123.590 1324.840 ;
        RECT 1124.430 1321.280 1136.470 1324.840 ;
        RECT 1137.310 1321.280 1146.130 1324.840 ;
        RECT 1146.970 1321.280 1155.790 1324.840 ;
        RECT 1156.630 1321.280 1165.450 1324.840 ;
        RECT 1166.290 1321.280 1175.110 1324.840 ;
        RECT 1175.950 1321.280 1187.990 1324.840 ;
        RECT 1188.830 1321.280 1197.650 1324.840 ;
        RECT 1198.490 1321.280 1207.310 1324.840 ;
        RECT 1208.150 1321.280 1216.970 1324.840 ;
        RECT 1217.810 1321.280 1226.630 1324.840 ;
        RECT 1227.470 1321.280 1239.510 1324.840 ;
        RECT 1240.350 1321.280 1249.170 1324.840 ;
        RECT 1250.010 1321.280 1258.830 1324.840 ;
        RECT 1259.670 1321.280 1268.490 1324.840 ;
        RECT 1269.330 1321.280 1278.150 1324.840 ;
        RECT 1278.990 1321.280 1291.030 1324.840 ;
        RECT 1291.870 1321.280 1300.690 1324.840 ;
        RECT 1301.530 1321.280 1310.350 1324.840 ;
        RECT 1311.190 1321.280 1314.580 1324.840 ;
        RECT 0.100 4.280 1314.580 1321.280 ;
        RECT 0.650 2.730 9.470 4.280 ;
        RECT 10.310 2.730 19.130 4.280 ;
        RECT 19.970 2.730 28.790 4.280 ;
        RECT 29.630 2.730 38.450 4.280 ;
        RECT 39.290 2.730 48.110 4.280 ;
        RECT 48.950 2.730 60.990 4.280 ;
        RECT 61.830 2.730 70.650 4.280 ;
        RECT 71.490 2.730 80.310 4.280 ;
        RECT 81.150 2.730 89.970 4.280 ;
        RECT 90.810 2.730 99.630 4.280 ;
        RECT 100.470 2.730 112.510 4.280 ;
        RECT 113.350 2.730 122.170 4.280 ;
        RECT 123.010 2.730 131.830 4.280 ;
        RECT 132.670 2.730 141.490 4.280 ;
        RECT 142.330 2.730 151.150 4.280 ;
        RECT 151.990 2.730 164.030 4.280 ;
        RECT 164.870 2.730 173.690 4.280 ;
        RECT 174.530 2.730 183.350 4.280 ;
        RECT 184.190 2.730 193.010 4.280 ;
        RECT 193.850 2.730 202.670 4.280 ;
        RECT 203.510 2.730 212.330 4.280 ;
        RECT 213.170 2.730 225.210 4.280 ;
        RECT 226.050 2.730 234.870 4.280 ;
        RECT 235.710 2.730 244.530 4.280 ;
        RECT 245.370 2.730 254.190 4.280 ;
        RECT 255.030 2.730 263.850 4.280 ;
        RECT 264.690 2.730 276.730 4.280 ;
        RECT 277.570 2.730 286.390 4.280 ;
        RECT 287.230 2.730 296.050 4.280 ;
        RECT 296.890 2.730 305.710 4.280 ;
        RECT 306.550 2.730 315.370 4.280 ;
        RECT 316.210 2.730 328.250 4.280 ;
        RECT 329.090 2.730 337.910 4.280 ;
        RECT 338.750 2.730 347.570 4.280 ;
        RECT 348.410 2.730 357.230 4.280 ;
        RECT 358.070 2.730 366.890 4.280 ;
        RECT 367.730 2.730 379.770 4.280 ;
        RECT 380.610 2.730 389.430 4.280 ;
        RECT 390.270 2.730 399.090 4.280 ;
        RECT 399.930 2.730 408.750 4.280 ;
        RECT 409.590 2.730 418.410 4.280 ;
        RECT 419.250 2.730 428.070 4.280 ;
        RECT 428.910 2.730 440.950 4.280 ;
        RECT 441.790 2.730 450.610 4.280 ;
        RECT 451.450 2.730 460.270 4.280 ;
        RECT 461.110 2.730 469.930 4.280 ;
        RECT 470.770 2.730 479.590 4.280 ;
        RECT 480.430 2.730 492.470 4.280 ;
        RECT 493.310 2.730 502.130 4.280 ;
        RECT 502.970 2.730 511.790 4.280 ;
        RECT 512.630 2.730 521.450 4.280 ;
        RECT 522.290 2.730 531.110 4.280 ;
        RECT 531.950 2.730 543.990 4.280 ;
        RECT 544.830 2.730 553.650 4.280 ;
        RECT 554.490 2.730 563.310 4.280 ;
        RECT 564.150 2.730 572.970 4.280 ;
        RECT 573.810 2.730 582.630 4.280 ;
        RECT 583.470 2.730 592.290 4.280 ;
        RECT 593.130 2.730 605.170 4.280 ;
        RECT 606.010 2.730 614.830 4.280 ;
        RECT 615.670 2.730 624.490 4.280 ;
        RECT 625.330 2.730 634.150 4.280 ;
        RECT 634.990 2.730 643.810 4.280 ;
        RECT 644.650 2.730 656.690 4.280 ;
        RECT 657.530 2.730 666.350 4.280 ;
        RECT 667.190 2.730 676.010 4.280 ;
        RECT 676.850 2.730 685.670 4.280 ;
        RECT 686.510 2.730 695.330 4.280 ;
        RECT 696.170 2.730 708.210 4.280 ;
        RECT 709.050 2.730 717.870 4.280 ;
        RECT 718.710 2.730 727.530 4.280 ;
        RECT 728.370 2.730 737.190 4.280 ;
        RECT 738.030 2.730 746.850 4.280 ;
        RECT 747.690 2.730 759.730 4.280 ;
        RECT 760.570 2.730 769.390 4.280 ;
        RECT 770.230 2.730 779.050 4.280 ;
        RECT 779.890 2.730 788.710 4.280 ;
        RECT 789.550 2.730 798.370 4.280 ;
        RECT 799.210 2.730 808.030 4.280 ;
        RECT 808.870 2.730 820.910 4.280 ;
        RECT 821.750 2.730 830.570 4.280 ;
        RECT 831.410 2.730 840.230 4.280 ;
        RECT 841.070 2.730 849.890 4.280 ;
        RECT 850.730 2.730 859.550 4.280 ;
        RECT 860.390 2.730 872.430 4.280 ;
        RECT 873.270 2.730 882.090 4.280 ;
        RECT 882.930 2.730 891.750 4.280 ;
        RECT 892.590 2.730 901.410 4.280 ;
        RECT 902.250 2.730 911.070 4.280 ;
        RECT 911.910 2.730 923.950 4.280 ;
        RECT 924.790 2.730 933.610 4.280 ;
        RECT 934.450 2.730 943.270 4.280 ;
        RECT 944.110 2.730 952.930 4.280 ;
        RECT 953.770 2.730 962.590 4.280 ;
        RECT 963.430 2.730 975.470 4.280 ;
        RECT 976.310 2.730 985.130 4.280 ;
        RECT 985.970 2.730 994.790 4.280 ;
        RECT 995.630 2.730 1004.450 4.280 ;
        RECT 1005.290 2.730 1014.110 4.280 ;
        RECT 1014.950 2.730 1023.770 4.280 ;
        RECT 1024.610 2.730 1036.650 4.280 ;
        RECT 1037.490 2.730 1046.310 4.280 ;
        RECT 1047.150 2.730 1055.970 4.280 ;
        RECT 1056.810 2.730 1065.630 4.280 ;
        RECT 1066.470 2.730 1075.290 4.280 ;
        RECT 1076.130 2.730 1088.170 4.280 ;
        RECT 1089.010 2.730 1097.830 4.280 ;
        RECT 1098.670 2.730 1107.490 4.280 ;
        RECT 1108.330 2.730 1117.150 4.280 ;
        RECT 1117.990 2.730 1126.810 4.280 ;
        RECT 1127.650 2.730 1139.690 4.280 ;
        RECT 1140.530 2.730 1149.350 4.280 ;
        RECT 1150.190 2.730 1159.010 4.280 ;
        RECT 1159.850 2.730 1168.670 4.280 ;
        RECT 1169.510 2.730 1178.330 4.280 ;
        RECT 1179.170 2.730 1187.990 4.280 ;
        RECT 1188.830 2.730 1200.870 4.280 ;
        RECT 1201.710 2.730 1210.530 4.280 ;
        RECT 1211.370 2.730 1220.190 4.280 ;
        RECT 1221.030 2.730 1229.850 4.280 ;
        RECT 1230.690 2.730 1239.510 4.280 ;
        RECT 1240.350 2.730 1252.390 4.280 ;
        RECT 1253.230 2.730 1262.050 4.280 ;
        RECT 1262.890 2.730 1271.710 4.280 ;
        RECT 1272.550 2.730 1281.370 4.280 ;
        RECT 1282.210 2.730 1291.030 4.280 ;
        RECT 1291.870 2.730 1303.910 4.280 ;
        RECT 1304.750 2.730 1313.570 4.280 ;
        RECT 1314.410 2.730 1314.580 4.280 ;
      LAYER met3 ;
        RECT 4.400 1322.240 1313.695 1323.105 ;
        RECT 3.950 1320.240 1313.695 1322.240 ;
        RECT 3.950 1318.840 1310.440 1320.240 ;
        RECT 3.950 1310.040 1313.695 1318.840 ;
        RECT 4.400 1308.640 1310.440 1310.040 ;
        RECT 3.950 1299.840 1313.695 1308.640 ;
        RECT 4.400 1298.440 1310.440 1299.840 ;
        RECT 3.950 1289.640 1313.695 1298.440 ;
        RECT 4.400 1288.240 1313.695 1289.640 ;
        RECT 3.950 1286.240 1313.695 1288.240 ;
        RECT 3.950 1284.840 1310.440 1286.240 ;
        RECT 3.950 1279.440 1313.695 1284.840 ;
        RECT 4.400 1278.040 1313.695 1279.440 ;
        RECT 3.950 1276.040 1313.695 1278.040 ;
        RECT 3.950 1274.640 1310.440 1276.040 ;
        RECT 3.950 1269.240 1313.695 1274.640 ;
        RECT 4.400 1267.840 1313.695 1269.240 ;
        RECT 3.950 1265.840 1313.695 1267.840 ;
        RECT 3.950 1264.440 1310.440 1265.840 ;
        RECT 3.950 1255.640 1313.695 1264.440 ;
        RECT 4.400 1254.240 1310.440 1255.640 ;
        RECT 3.950 1245.440 1313.695 1254.240 ;
        RECT 4.400 1244.040 1310.440 1245.440 ;
        RECT 3.950 1235.240 1313.695 1244.040 ;
        RECT 4.400 1233.840 1313.695 1235.240 ;
        RECT 3.950 1231.840 1313.695 1233.840 ;
        RECT 3.950 1230.440 1310.440 1231.840 ;
        RECT 3.950 1225.040 1313.695 1230.440 ;
        RECT 4.400 1223.640 1313.695 1225.040 ;
        RECT 3.950 1221.640 1313.695 1223.640 ;
        RECT 3.950 1220.240 1310.440 1221.640 ;
        RECT 3.950 1214.840 1313.695 1220.240 ;
        RECT 4.400 1213.440 1313.695 1214.840 ;
        RECT 3.950 1211.440 1313.695 1213.440 ;
        RECT 3.950 1210.040 1310.440 1211.440 ;
        RECT 3.950 1204.640 1313.695 1210.040 ;
        RECT 4.400 1203.240 1313.695 1204.640 ;
        RECT 3.950 1201.240 1313.695 1203.240 ;
        RECT 3.950 1199.840 1310.440 1201.240 ;
        RECT 3.950 1191.040 1313.695 1199.840 ;
        RECT 4.400 1189.640 1310.440 1191.040 ;
        RECT 3.950 1180.840 1313.695 1189.640 ;
        RECT 4.400 1179.440 1313.695 1180.840 ;
        RECT 3.950 1177.440 1313.695 1179.440 ;
        RECT 3.950 1176.040 1310.440 1177.440 ;
        RECT 3.950 1170.640 1313.695 1176.040 ;
        RECT 4.400 1169.240 1313.695 1170.640 ;
        RECT 3.950 1167.240 1313.695 1169.240 ;
        RECT 3.950 1165.840 1310.440 1167.240 ;
        RECT 3.950 1160.440 1313.695 1165.840 ;
        RECT 4.400 1159.040 1313.695 1160.440 ;
        RECT 3.950 1157.040 1313.695 1159.040 ;
        RECT 3.950 1155.640 1310.440 1157.040 ;
        RECT 3.950 1150.240 1313.695 1155.640 ;
        RECT 4.400 1148.840 1313.695 1150.240 ;
        RECT 3.950 1146.840 1313.695 1148.840 ;
        RECT 3.950 1145.440 1310.440 1146.840 ;
        RECT 3.950 1136.640 1313.695 1145.440 ;
        RECT 4.400 1135.240 1310.440 1136.640 ;
        RECT 3.950 1126.440 1313.695 1135.240 ;
        RECT 4.400 1125.040 1313.695 1126.440 ;
        RECT 3.950 1123.040 1313.695 1125.040 ;
        RECT 3.950 1121.640 1310.440 1123.040 ;
        RECT 3.950 1116.240 1313.695 1121.640 ;
        RECT 4.400 1114.840 1313.695 1116.240 ;
        RECT 3.950 1112.840 1313.695 1114.840 ;
        RECT 3.950 1111.440 1310.440 1112.840 ;
        RECT 3.950 1106.040 1313.695 1111.440 ;
        RECT 4.400 1104.640 1313.695 1106.040 ;
        RECT 3.950 1102.640 1313.695 1104.640 ;
        RECT 3.950 1101.240 1310.440 1102.640 ;
        RECT 3.950 1095.840 1313.695 1101.240 ;
        RECT 4.400 1094.440 1313.695 1095.840 ;
        RECT 3.950 1092.440 1313.695 1094.440 ;
        RECT 3.950 1091.040 1310.440 1092.440 ;
        RECT 3.950 1082.240 1313.695 1091.040 ;
        RECT 4.400 1080.840 1310.440 1082.240 ;
        RECT 3.950 1072.040 1313.695 1080.840 ;
        RECT 4.400 1070.640 1310.440 1072.040 ;
        RECT 3.950 1061.840 1313.695 1070.640 ;
        RECT 4.400 1060.440 1313.695 1061.840 ;
        RECT 3.950 1058.440 1313.695 1060.440 ;
        RECT 3.950 1057.040 1310.440 1058.440 ;
        RECT 3.950 1051.640 1313.695 1057.040 ;
        RECT 4.400 1050.240 1313.695 1051.640 ;
        RECT 3.950 1048.240 1313.695 1050.240 ;
        RECT 3.950 1046.840 1310.440 1048.240 ;
        RECT 3.950 1041.440 1313.695 1046.840 ;
        RECT 4.400 1040.040 1313.695 1041.440 ;
        RECT 3.950 1038.040 1313.695 1040.040 ;
        RECT 3.950 1036.640 1310.440 1038.040 ;
        RECT 3.950 1031.240 1313.695 1036.640 ;
        RECT 4.400 1029.840 1313.695 1031.240 ;
        RECT 3.950 1027.840 1313.695 1029.840 ;
        RECT 3.950 1026.440 1310.440 1027.840 ;
        RECT 3.950 1017.640 1313.695 1026.440 ;
        RECT 4.400 1016.240 1310.440 1017.640 ;
        RECT 3.950 1007.440 1313.695 1016.240 ;
        RECT 4.400 1006.040 1313.695 1007.440 ;
        RECT 3.950 1004.040 1313.695 1006.040 ;
        RECT 3.950 1002.640 1310.440 1004.040 ;
        RECT 3.950 997.240 1313.695 1002.640 ;
        RECT 4.400 995.840 1313.695 997.240 ;
        RECT 3.950 993.840 1313.695 995.840 ;
        RECT 3.950 992.440 1310.440 993.840 ;
        RECT 3.950 987.040 1313.695 992.440 ;
        RECT 4.400 985.640 1313.695 987.040 ;
        RECT 3.950 983.640 1313.695 985.640 ;
        RECT 3.950 982.240 1310.440 983.640 ;
        RECT 3.950 976.840 1313.695 982.240 ;
        RECT 4.400 975.440 1313.695 976.840 ;
        RECT 3.950 973.440 1313.695 975.440 ;
        RECT 3.950 972.040 1310.440 973.440 ;
        RECT 3.950 963.240 1313.695 972.040 ;
        RECT 4.400 961.840 1310.440 963.240 ;
        RECT 3.950 953.040 1313.695 961.840 ;
        RECT 4.400 951.640 1313.695 953.040 ;
        RECT 3.950 949.640 1313.695 951.640 ;
        RECT 3.950 948.240 1310.440 949.640 ;
        RECT 3.950 942.840 1313.695 948.240 ;
        RECT 4.400 941.440 1313.695 942.840 ;
        RECT 3.950 939.440 1313.695 941.440 ;
        RECT 3.950 938.040 1310.440 939.440 ;
        RECT 3.950 932.640 1313.695 938.040 ;
        RECT 4.400 931.240 1313.695 932.640 ;
        RECT 3.950 929.240 1313.695 931.240 ;
        RECT 3.950 927.840 1310.440 929.240 ;
        RECT 3.950 922.440 1313.695 927.840 ;
        RECT 4.400 921.040 1313.695 922.440 ;
        RECT 3.950 919.040 1313.695 921.040 ;
        RECT 3.950 917.640 1310.440 919.040 ;
        RECT 3.950 908.840 1313.695 917.640 ;
        RECT 4.400 907.440 1310.440 908.840 ;
        RECT 3.950 898.640 1313.695 907.440 ;
        RECT 4.400 897.240 1310.440 898.640 ;
        RECT 3.950 888.440 1313.695 897.240 ;
        RECT 4.400 887.040 1313.695 888.440 ;
        RECT 3.950 885.040 1313.695 887.040 ;
        RECT 3.950 883.640 1310.440 885.040 ;
        RECT 3.950 878.240 1313.695 883.640 ;
        RECT 4.400 876.840 1313.695 878.240 ;
        RECT 3.950 874.840 1313.695 876.840 ;
        RECT 3.950 873.440 1310.440 874.840 ;
        RECT 3.950 868.040 1313.695 873.440 ;
        RECT 4.400 866.640 1313.695 868.040 ;
        RECT 3.950 864.640 1313.695 866.640 ;
        RECT 3.950 863.240 1310.440 864.640 ;
        RECT 3.950 854.440 1313.695 863.240 ;
        RECT 4.400 853.040 1310.440 854.440 ;
        RECT 3.950 844.240 1313.695 853.040 ;
        RECT 4.400 842.840 1310.440 844.240 ;
        RECT 3.950 834.040 1313.695 842.840 ;
        RECT 4.400 832.640 1313.695 834.040 ;
        RECT 3.950 830.640 1313.695 832.640 ;
        RECT 3.950 829.240 1310.440 830.640 ;
        RECT 3.950 823.840 1313.695 829.240 ;
        RECT 4.400 822.440 1313.695 823.840 ;
        RECT 3.950 820.440 1313.695 822.440 ;
        RECT 3.950 819.040 1310.440 820.440 ;
        RECT 3.950 813.640 1313.695 819.040 ;
        RECT 4.400 812.240 1313.695 813.640 ;
        RECT 3.950 810.240 1313.695 812.240 ;
        RECT 3.950 808.840 1310.440 810.240 ;
        RECT 3.950 803.440 1313.695 808.840 ;
        RECT 4.400 802.040 1313.695 803.440 ;
        RECT 3.950 800.040 1313.695 802.040 ;
        RECT 3.950 798.640 1310.440 800.040 ;
        RECT 3.950 789.840 1313.695 798.640 ;
        RECT 4.400 788.440 1310.440 789.840 ;
        RECT 3.950 779.640 1313.695 788.440 ;
        RECT 4.400 778.240 1313.695 779.640 ;
        RECT 3.950 776.240 1313.695 778.240 ;
        RECT 3.950 774.840 1310.440 776.240 ;
        RECT 3.950 769.440 1313.695 774.840 ;
        RECT 4.400 768.040 1313.695 769.440 ;
        RECT 3.950 766.040 1313.695 768.040 ;
        RECT 3.950 764.640 1310.440 766.040 ;
        RECT 3.950 759.240 1313.695 764.640 ;
        RECT 4.400 757.840 1313.695 759.240 ;
        RECT 3.950 755.840 1313.695 757.840 ;
        RECT 3.950 754.440 1310.440 755.840 ;
        RECT 3.950 749.040 1313.695 754.440 ;
        RECT 4.400 747.640 1313.695 749.040 ;
        RECT 3.950 745.640 1313.695 747.640 ;
        RECT 3.950 744.240 1310.440 745.640 ;
        RECT 3.950 735.440 1313.695 744.240 ;
        RECT 4.400 734.040 1310.440 735.440 ;
        RECT 3.950 725.240 1313.695 734.040 ;
        RECT 4.400 723.840 1313.695 725.240 ;
        RECT 3.950 721.840 1313.695 723.840 ;
        RECT 3.950 720.440 1310.440 721.840 ;
        RECT 3.950 715.040 1313.695 720.440 ;
        RECT 4.400 713.640 1313.695 715.040 ;
        RECT 3.950 711.640 1313.695 713.640 ;
        RECT 3.950 710.240 1310.440 711.640 ;
        RECT 3.950 704.840 1313.695 710.240 ;
        RECT 4.400 703.440 1313.695 704.840 ;
        RECT 3.950 701.440 1313.695 703.440 ;
        RECT 3.950 700.040 1310.440 701.440 ;
        RECT 3.950 694.640 1313.695 700.040 ;
        RECT 4.400 693.240 1313.695 694.640 ;
        RECT 3.950 691.240 1313.695 693.240 ;
        RECT 3.950 689.840 1310.440 691.240 ;
        RECT 3.950 681.040 1313.695 689.840 ;
        RECT 4.400 679.640 1310.440 681.040 ;
        RECT 3.950 670.840 1313.695 679.640 ;
        RECT 4.400 669.440 1310.440 670.840 ;
        RECT 3.950 660.640 1313.695 669.440 ;
        RECT 4.400 659.240 1313.695 660.640 ;
        RECT 3.950 657.240 1313.695 659.240 ;
        RECT 3.950 655.840 1310.440 657.240 ;
        RECT 3.950 650.440 1313.695 655.840 ;
        RECT 4.400 649.040 1313.695 650.440 ;
        RECT 3.950 647.040 1313.695 649.040 ;
        RECT 3.950 645.640 1310.440 647.040 ;
        RECT 3.950 640.240 1313.695 645.640 ;
        RECT 4.400 638.840 1313.695 640.240 ;
        RECT 3.950 636.840 1313.695 638.840 ;
        RECT 3.950 635.440 1310.440 636.840 ;
        RECT 3.950 626.640 1313.695 635.440 ;
        RECT 4.400 625.240 1310.440 626.640 ;
        RECT 3.950 616.440 1313.695 625.240 ;
        RECT 4.400 615.040 1310.440 616.440 ;
        RECT 3.950 606.240 1313.695 615.040 ;
        RECT 4.400 604.840 1313.695 606.240 ;
        RECT 3.950 602.840 1313.695 604.840 ;
        RECT 3.950 601.440 1310.440 602.840 ;
        RECT 3.950 596.040 1313.695 601.440 ;
        RECT 4.400 594.640 1313.695 596.040 ;
        RECT 3.950 592.640 1313.695 594.640 ;
        RECT 3.950 591.240 1310.440 592.640 ;
        RECT 3.950 585.840 1313.695 591.240 ;
        RECT 4.400 584.440 1313.695 585.840 ;
        RECT 3.950 582.440 1313.695 584.440 ;
        RECT 3.950 581.040 1310.440 582.440 ;
        RECT 3.950 575.640 1313.695 581.040 ;
        RECT 4.400 574.240 1313.695 575.640 ;
        RECT 3.950 572.240 1313.695 574.240 ;
        RECT 3.950 570.840 1310.440 572.240 ;
        RECT 3.950 562.040 1313.695 570.840 ;
        RECT 4.400 560.640 1310.440 562.040 ;
        RECT 3.950 551.840 1313.695 560.640 ;
        RECT 4.400 550.440 1313.695 551.840 ;
        RECT 3.950 548.440 1313.695 550.440 ;
        RECT 3.950 547.040 1310.440 548.440 ;
        RECT 3.950 541.640 1313.695 547.040 ;
        RECT 4.400 540.240 1313.695 541.640 ;
        RECT 3.950 538.240 1313.695 540.240 ;
        RECT 3.950 536.840 1310.440 538.240 ;
        RECT 3.950 531.440 1313.695 536.840 ;
        RECT 4.400 530.040 1313.695 531.440 ;
        RECT 3.950 528.040 1313.695 530.040 ;
        RECT 3.950 526.640 1310.440 528.040 ;
        RECT 3.950 521.240 1313.695 526.640 ;
        RECT 4.400 519.840 1313.695 521.240 ;
        RECT 3.950 517.840 1313.695 519.840 ;
        RECT 3.950 516.440 1310.440 517.840 ;
        RECT 3.950 507.640 1313.695 516.440 ;
        RECT 4.400 506.240 1310.440 507.640 ;
        RECT 3.950 497.440 1313.695 506.240 ;
        RECT 4.400 496.040 1313.695 497.440 ;
        RECT 3.950 494.040 1313.695 496.040 ;
        RECT 3.950 492.640 1310.440 494.040 ;
        RECT 3.950 487.240 1313.695 492.640 ;
        RECT 4.400 485.840 1313.695 487.240 ;
        RECT 3.950 483.840 1313.695 485.840 ;
        RECT 3.950 482.440 1310.440 483.840 ;
        RECT 3.950 477.040 1313.695 482.440 ;
        RECT 4.400 475.640 1313.695 477.040 ;
        RECT 3.950 473.640 1313.695 475.640 ;
        RECT 3.950 472.240 1310.440 473.640 ;
        RECT 3.950 466.840 1313.695 472.240 ;
        RECT 4.400 465.440 1313.695 466.840 ;
        RECT 3.950 463.440 1313.695 465.440 ;
        RECT 3.950 462.040 1310.440 463.440 ;
        RECT 3.950 453.240 1313.695 462.040 ;
        RECT 4.400 451.840 1310.440 453.240 ;
        RECT 3.950 443.040 1313.695 451.840 ;
        RECT 4.400 441.640 1310.440 443.040 ;
        RECT 3.950 432.840 1313.695 441.640 ;
        RECT 4.400 431.440 1313.695 432.840 ;
        RECT 3.950 429.440 1313.695 431.440 ;
        RECT 3.950 428.040 1310.440 429.440 ;
        RECT 3.950 422.640 1313.695 428.040 ;
        RECT 4.400 421.240 1313.695 422.640 ;
        RECT 3.950 419.240 1313.695 421.240 ;
        RECT 3.950 417.840 1310.440 419.240 ;
        RECT 3.950 412.440 1313.695 417.840 ;
        RECT 4.400 411.040 1313.695 412.440 ;
        RECT 3.950 409.040 1313.695 411.040 ;
        RECT 3.950 407.640 1310.440 409.040 ;
        RECT 3.950 402.240 1313.695 407.640 ;
        RECT 4.400 400.840 1313.695 402.240 ;
        RECT 3.950 398.840 1313.695 400.840 ;
        RECT 3.950 397.440 1310.440 398.840 ;
        RECT 3.950 388.640 1313.695 397.440 ;
        RECT 4.400 387.240 1310.440 388.640 ;
        RECT 3.950 378.440 1313.695 387.240 ;
        RECT 4.400 377.040 1313.695 378.440 ;
        RECT 3.950 375.040 1313.695 377.040 ;
        RECT 3.950 373.640 1310.440 375.040 ;
        RECT 3.950 368.240 1313.695 373.640 ;
        RECT 4.400 366.840 1313.695 368.240 ;
        RECT 3.950 364.840 1313.695 366.840 ;
        RECT 3.950 363.440 1310.440 364.840 ;
        RECT 3.950 358.040 1313.695 363.440 ;
        RECT 4.400 356.640 1313.695 358.040 ;
        RECT 3.950 354.640 1313.695 356.640 ;
        RECT 3.950 353.240 1310.440 354.640 ;
        RECT 3.950 347.840 1313.695 353.240 ;
        RECT 4.400 346.440 1313.695 347.840 ;
        RECT 3.950 344.440 1313.695 346.440 ;
        RECT 3.950 343.040 1310.440 344.440 ;
        RECT 3.950 334.240 1313.695 343.040 ;
        RECT 4.400 332.840 1310.440 334.240 ;
        RECT 3.950 324.040 1313.695 332.840 ;
        RECT 4.400 322.640 1313.695 324.040 ;
        RECT 3.950 320.640 1313.695 322.640 ;
        RECT 3.950 319.240 1310.440 320.640 ;
        RECT 3.950 313.840 1313.695 319.240 ;
        RECT 4.400 312.440 1313.695 313.840 ;
        RECT 3.950 310.440 1313.695 312.440 ;
        RECT 3.950 309.040 1310.440 310.440 ;
        RECT 3.950 303.640 1313.695 309.040 ;
        RECT 4.400 302.240 1313.695 303.640 ;
        RECT 3.950 300.240 1313.695 302.240 ;
        RECT 3.950 298.840 1310.440 300.240 ;
        RECT 3.950 293.440 1313.695 298.840 ;
        RECT 4.400 292.040 1313.695 293.440 ;
        RECT 3.950 290.040 1313.695 292.040 ;
        RECT 3.950 288.640 1310.440 290.040 ;
        RECT 3.950 279.840 1313.695 288.640 ;
        RECT 4.400 278.440 1310.440 279.840 ;
        RECT 3.950 269.640 1313.695 278.440 ;
        RECT 4.400 268.240 1310.440 269.640 ;
        RECT 3.950 259.440 1313.695 268.240 ;
        RECT 4.400 258.040 1313.695 259.440 ;
        RECT 3.950 256.040 1313.695 258.040 ;
        RECT 3.950 254.640 1310.440 256.040 ;
        RECT 3.950 249.240 1313.695 254.640 ;
        RECT 4.400 247.840 1313.695 249.240 ;
        RECT 3.950 245.840 1313.695 247.840 ;
        RECT 3.950 244.440 1310.440 245.840 ;
        RECT 3.950 239.040 1313.695 244.440 ;
        RECT 4.400 237.640 1313.695 239.040 ;
        RECT 3.950 235.640 1313.695 237.640 ;
        RECT 3.950 234.240 1310.440 235.640 ;
        RECT 3.950 225.440 1313.695 234.240 ;
        RECT 4.400 224.040 1310.440 225.440 ;
        RECT 3.950 215.240 1313.695 224.040 ;
        RECT 4.400 213.840 1310.440 215.240 ;
        RECT 3.950 205.040 1313.695 213.840 ;
        RECT 4.400 203.640 1313.695 205.040 ;
        RECT 3.950 201.640 1313.695 203.640 ;
        RECT 3.950 200.240 1310.440 201.640 ;
        RECT 3.950 194.840 1313.695 200.240 ;
        RECT 4.400 193.440 1313.695 194.840 ;
        RECT 3.950 191.440 1313.695 193.440 ;
        RECT 3.950 190.040 1310.440 191.440 ;
        RECT 3.950 184.640 1313.695 190.040 ;
        RECT 4.400 183.240 1313.695 184.640 ;
        RECT 3.950 181.240 1313.695 183.240 ;
        RECT 3.950 179.840 1310.440 181.240 ;
        RECT 3.950 174.440 1313.695 179.840 ;
        RECT 4.400 173.040 1313.695 174.440 ;
        RECT 3.950 171.040 1313.695 173.040 ;
        RECT 3.950 169.640 1310.440 171.040 ;
        RECT 3.950 160.840 1313.695 169.640 ;
        RECT 4.400 159.440 1310.440 160.840 ;
        RECT 3.950 150.640 1313.695 159.440 ;
        RECT 4.400 149.240 1313.695 150.640 ;
        RECT 3.950 147.240 1313.695 149.240 ;
        RECT 3.950 145.840 1310.440 147.240 ;
        RECT 3.950 140.440 1313.695 145.840 ;
        RECT 4.400 139.040 1313.695 140.440 ;
        RECT 3.950 137.040 1313.695 139.040 ;
        RECT 3.950 135.640 1310.440 137.040 ;
        RECT 3.950 130.240 1313.695 135.640 ;
        RECT 4.400 128.840 1313.695 130.240 ;
        RECT 3.950 126.840 1313.695 128.840 ;
        RECT 3.950 125.440 1310.440 126.840 ;
        RECT 3.950 120.040 1313.695 125.440 ;
        RECT 4.400 118.640 1313.695 120.040 ;
        RECT 3.950 116.640 1313.695 118.640 ;
        RECT 3.950 115.240 1310.440 116.640 ;
        RECT 3.950 106.440 1313.695 115.240 ;
        RECT 4.400 105.040 1310.440 106.440 ;
        RECT 3.950 96.240 1313.695 105.040 ;
        RECT 4.400 94.840 1313.695 96.240 ;
        RECT 3.950 92.840 1313.695 94.840 ;
        RECT 3.950 91.440 1310.440 92.840 ;
        RECT 3.950 86.040 1313.695 91.440 ;
        RECT 4.400 84.640 1313.695 86.040 ;
        RECT 3.950 82.640 1313.695 84.640 ;
        RECT 3.950 81.240 1310.440 82.640 ;
        RECT 3.950 75.840 1313.695 81.240 ;
        RECT 4.400 74.440 1313.695 75.840 ;
        RECT 3.950 72.440 1313.695 74.440 ;
        RECT 3.950 71.040 1310.440 72.440 ;
        RECT 3.950 65.640 1313.695 71.040 ;
        RECT 4.400 64.240 1313.695 65.640 ;
        RECT 3.950 62.240 1313.695 64.240 ;
        RECT 3.950 60.840 1310.440 62.240 ;
        RECT 3.950 52.040 1313.695 60.840 ;
        RECT 4.400 50.640 1310.440 52.040 ;
        RECT 3.950 41.840 1313.695 50.640 ;
        RECT 4.400 40.440 1310.440 41.840 ;
        RECT 3.950 31.640 1313.695 40.440 ;
        RECT 4.400 30.240 1313.695 31.640 ;
        RECT 3.950 28.240 1313.695 30.240 ;
        RECT 3.950 26.840 1310.440 28.240 ;
        RECT 3.950 21.440 1313.695 26.840 ;
        RECT 4.400 20.040 1313.695 21.440 ;
        RECT 3.950 18.040 1313.695 20.040 ;
        RECT 3.950 16.640 1310.440 18.040 ;
        RECT 3.950 11.240 1313.695 16.640 ;
        RECT 4.400 9.840 1313.695 11.240 ;
        RECT 3.950 7.840 1313.695 9.840 ;
        RECT 3.950 6.440 1310.440 7.840 ;
        RECT 3.950 6.295 1313.695 6.440 ;
      LAYER met4 ;
        RECT 3.550 1314.400 1303.345 1316.985 ;
        RECT 3.550 10.240 20.640 1314.400 ;
        RECT 23.040 10.240 23.940 1314.400 ;
        RECT 26.340 10.240 174.240 1314.400 ;
        RECT 176.640 10.240 177.540 1314.400 ;
        RECT 179.940 10.240 327.840 1314.400 ;
        RECT 330.240 10.240 331.140 1314.400 ;
        RECT 333.540 10.240 481.440 1314.400 ;
        RECT 483.840 10.240 484.740 1314.400 ;
        RECT 487.140 10.240 635.040 1314.400 ;
        RECT 637.440 10.240 638.340 1314.400 ;
        RECT 640.740 10.240 788.640 1314.400 ;
        RECT 791.040 10.240 791.940 1314.400 ;
        RECT 794.340 10.240 942.240 1314.400 ;
        RECT 944.640 10.240 945.540 1314.400 ;
        RECT 947.940 10.240 1095.840 1314.400 ;
        RECT 1098.240 10.240 1099.140 1314.400 ;
        RECT 1101.540 10.240 1249.440 1314.400 ;
        RECT 1251.840 10.240 1252.740 1314.400 ;
        RECT 1255.140 10.240 1303.345 1314.400 ;
        RECT 3.550 6.295 1303.345 10.240 ;
      LAYER met5 ;
        RECT 3.340 799.130 1287.420 920.500 ;
        RECT 3.340 791.030 3.680 799.130 ;
        RECT 3.340 645.950 1287.420 791.030 ;
        RECT 3.340 637.850 3.680 645.950 ;
        RECT 3.340 492.770 1287.420 637.850 ;
        RECT 3.340 484.670 3.680 492.770 ;
        RECT 3.340 339.590 1287.420 484.670 ;
        RECT 3.340 331.490 3.680 339.590 ;
        RECT 3.340 186.410 1287.420 331.490 ;
        RECT 3.340 178.310 3.680 186.410 ;
        RECT 3.340 174.300 1287.420 178.310 ;
  END
END D2DAdapter
END LIBRARY

